// Register File:
module RegisterFile
(
	
);

endmodule