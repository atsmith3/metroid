module Bit_Serial_Processor(input [1:0] R,
									 input Execute, LoadA, LoadB, Reset, Clk,
									 input [2:0] F,
									 output [7:0] Aval, Bval,
									 output [6:0] AhexU, AhexL, BhexU, BhexL,
									 output [3:0] LED);
				testbench_8	test0();
endmodule