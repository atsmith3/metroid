// Controller logic 8 bit multiplier

module Controller(	input logic ClearA_LoadB, Run, Reset, Clk,
							output logic Clr_Ld, Load, Shift, Add, Sub);
							

							
endmodule


