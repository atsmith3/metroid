module kraid(
	input logic  			kraid_r_en, kraid_g_en, kraid_n_en, kraid_shoot_en, kraid_throw_en, kraid_throw_2_en, kraid_dir, kraid_as_dir,
	input logic  [10:0] 	vga_x, vga_y, kraid_y, kraid_x, shoot_x, shoot_y, throw_x, throw_y, throw_2_x, throw_2_y,
	output logic [6:0] 	color,
	output logic 			draw
);

   parameter kraid_h = 62;
	parameter kraid_w = 46;
	
	parameter shoot_h = 18;
	parameter shoot_w = 21;
	
	parameter attack_h = 12;
	parameter attack_w = 17;

	logic [6:0] kraid_n[kraid_h][kraid_w];
	logic [6:0] kraid_r[kraid_h][kraid_w];
	logic [6:0] kraid_g[kraid_h][kraid_w];
	logic [6:0] shoot[shoot_h][shoot_w];
	logic [6:0] attack[attack_h][attack_w];
	
	always_ff begin
		kraid_r = '{'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,33,10,8,8,8,8,10,33,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,30,33,8,8,8,30,32,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,8,8,8,30,32,8,8,8,32,30,8,8,30,27,28,28,28,28,28,8,8,28,8,8,8,28,8,8,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,8,8,8,32,32,8,8,8,32,30,8,8,30,19,24,24,24,24,27,8,8,8,8,8,33,27,8,8,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,30,33,8,32,30,28,27,19,12,12,30,30,22,30,19,32,33,1,12,12,19,8,8,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,8,8,33,33,32,33,8,8,1,12,30,24,30,30,30,13,1,19,30,30,22,1,19,12,10,33,33,33,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,8,10,12,12,30,33,33,27,10,12,12,12,30,30,30,1,33,13,30,30,30,30,30,12,33,33,19,30,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,10,1,32,27,24,24,32,33,33,30,30,30,30,30,12,19,33,33,27,33,33,33,1,30,30,30,19,19,33,8,10,33,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,19,12,15,24,27,27,27,33,1,12,30,30,30,30,12,10,33,33,27,33,33,33,33,30,30,30,30,22,33,33,19,32,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,19,24,27,33,33,33,33,19,30,30,33,33,33,33,22,30,19,1,33,20,12,30,30,33,1,22,30,30,12,12,30,32,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,33,10,24,32,33,33,33,33,30,19,13,1,33,33,33,19,19,30,1,33,30,30,30,20,33,1,20,19,30,12,30,10,33,8,8,8,8,8,8},
						'{8,8,8,28,8,8,19,32,27,33,33,33,33,33,33,30,1,33,13,12,12,30,33,1,30,30,12,33,33,27,33,33,33,33,13,22,12,30,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,27,24,27,33,33,33,1,1,33,33,33,1,19,12,30,1,1,13,30,30,12,1,1,33,33,33,33,33,13,30,30,30,8,8,8,8,8,8,8,8},
						'{8,8,8,8,28,28,28,28,27,27,27,30,12,12,32,8,33,30,30,30,33,33,30,30,30,30,30,30,30,33,33,33,33,27,10,30,30,10,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,8,33,24,24,24,24,33,8,33,19,30,30,33,33,1,33,1,33,1,19,30,13,13,13,10,27,30,30,30,30,32,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,8,33,19,27,28,28,28,8,33,30,30,19,33,33,33,33,33,33,33,32,30,30,30,30,30,30,30,30,30,30,12,32,8,8,8,8,8,8},
						'{8,8,8,8,10,27,30,33,8,8,8,28,28,8,8,8,8,8,32,30,19,13,33,33,33,1,27,8,8,30,30,30,30,12,30,30,12,12,12,32,8,8,8,8,8,8},
						'{8,8,8,8,32,30,12,32,8,8,8,8,28,8,8,8,8,8,33,30,30,19,33,33,33,13,19,8,8,10,30,30,30,12,30,30,30,12,12,32,8,8,8,8,8,8},
						'{8,8,32,19,27,27,27,27,30,33,8,8,8,8,8,8,8,8,8,8,10,30,19,19,30,22,30,8,8,8,8,30,30,30,12,12,30,30,30,30,19,33,8,8,8,8},
						'{8,8,33,30,27,27,27,24,24,8,8,8,8,8,8,8,8,8,8,8,33,32,32,32,32,32,32,33,8,8,8,32,10,30,30,12,13,13,30,30,30,33,8,8,8,8},
						'{8,8,8,24,27,24,27,27,27,27,27,28,27,8,8,30,33,8,8,8,8,8,8,8,8,8,8,32,30,8,8,8,33,22,30,30,33,33,30,30,30,33,8,8,8,8},
						'{8,33,33,24,27,27,27,28,8,8,8,8,8,8,8,30,10,33,33,33,32,33,33,33,8,8,8,33,33,33,33,8,33,30,30,30,13,1,30,30,30,33,8,8,8,8},
						'{33,19,24,27,27,24,27,8,8,8,8,8,8,8,8,19,12,12,30,30,12,12,30,32,8,8,8,8,8,30,32,8,33,19,30,30,30,30,30,30,30,33,8,8,8,8},
						'{33,24,27,24,33,33,10,33,8,8,8,8,8,10,10,30,30,30,30,30,30,30,30,30,32,32,32,32,10,8,8,8,8,8,8,8,30,30,30,32,8,8,8,8,8,8},
						'{33,24,27,27,33,33,30,32,8,8,8,8,8,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,8,8,8,8,8,8,8,10,30,30,32,8,8,8,8,8,8},
						'{33,33,33,24,19,30,12,32,28,28,28,8,8,8,8,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,19,8,8,8,8,8,8,8,8,8,8,8,8},
						'{33,33,33,27,22,30,30,24,27,27,28,8,8,8,8,30,30,30,30,30,30,30,30,19,19,13,19,19,30,30,30,30,30,19,33,8,8,8,8,8,8,8,8,8,8,8},
						'{33,33,33,33,19,30,27,27,27,24,28,8,8,30,30,30,30,30,30,30,30,30,12,30,33,33,33,13,30,30,30,30,30,30,30,19,30,30,8,8,8,8,8,8,8,8},
						'{33,33,33,1,30,24,27,27,27,28,8,8,8,33,32,30,30,30,30,30,13,1,13,33,33,33,1,19,30,30,30,30,30,30,30,19,32,33,8,8,8,8,8,8,8,8},
						'{33,33,13,12,27,27,27,27,28,8,8,8,8,8,8,30,19,30,30,12,33,33,33,33,33,1,30,30,30,30,30,30,30,30,30,30,8,8,8,8,8,8,8,8,8,8},
						'{33,13,24,24,24,27,27,28,8,8,8,33,32,8,8,30,30,30,30,30,10,13,33,33,33,33,1,33,1,30,30,30,19,30,1,33,32,33,8,8,8,8,8,8,8,8},
						'{1,12,24,28,28,27,28,8,8,8,8,32,30,8,8,30,30,30,30,30,12,30,33,33,33,33,33,33,33,19,30,30,30,30,33,33,19,10,8,8,8,8,8,8,8,8},
						'{8,28,24,28,8,8,8,8,8,33,10,33,8,10,32,8,33,30,30,30,30,22,19,19,19,19,19,33,33,33,33,33,33,33,1,19,19,30,10,33,8,8,8,8,8,8},
						'{8,28,28,28,8,8,8,8,8,33,10,8,33,30,10,8,33,30,10,30,30,30,30,19,19,30,30,33,33,33,33,33,33,33,13,19,30,30,30,32,8,8,8,8,8,8},
						'{8,8,8,27,27,27,28,8,8,8,8,32,30,19,10,8,8,8,8,8,8,8,30,13,33,33,33,13,30,19,19,33,33,33,13,30,30,30,30,30,19,33,8,8,8,8},
						'{8,8,33,24,10,10,27,8,8,8,8,33,32,32,33,8,8,8,8,8,8,8,32,33,33,33,33,19,30,13,1,1,33,33,1,13,13,13,13,19,12,33,8,8,8,8},
						'{8,8,32,19,24,27,27,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,12,24,24,10,30,33,33,12,32,33,33,33,33,33,33,33,12,33,8,8,8,8},
						'{8,8,8,24,27,27,33,8,8,8,8,33,33,33,33,33,33,33,33,33,8,8,33,32,24,32,33,33,1,1,10,10,28,33,33,1,1,1,33,33,12,33,8,8,8,8},
						'{8,8,8,28,28,27,33,33,27,8,8,32,30,30,30,30,30,30,30,30,8,8,19,30,27,33,33,33,33,30,30,27,33,33,13,30,30,19,33,8,19,33,8,8,8,8},
						'{8,8,8,8,28,27,30,19,10,32,10,30,30,33,33,33,33,33,13,30,10,32,8,33,33,33,33,1,19,24,32,33,28,13,19,30,30,19,13,32,8,8,8,8,8,8},
						'{8,8,8,8,28,24,15,12,12,12,12,30,30,33,33,33,33,33,13,30,19,19,33,33,33,33,33,19,30,24,27,33,1,30,30,30,30,30,30,32,8,8,8,8,8,8},
						'{8,8,8,28,8,33,12,30,27,27,27,27,27,33,33,19,1,33,33,33,19,30,19,19,19,19,30,33,33,33,33,19,30,30,30,19,30,30,30,30,30,33,8,8,8,8},
						'{8,8,8,28,8,33,30,24,27,27,27,32,27,33,1,30,13,33,33,33,19,30,30,19,19,19,13,33,33,33,33,30,30,30,30,30,30,19,30,30,10,33,8,8,8,8},
						'{8,8,8,8,28,27,27,27,27,33,33,33,33,30,30,30,30,30,30,30,30,30,30,13,33,33,33,33,33,33,33,12,12,12,30,30,30,30,30,32,8,8,8,8,8,8},
						'{8,8,8,8,8,8,27,27,33,33,33,33,1,30,30,30,30,30,30,30,13,1,30,19,1,1,1,33,33,1,32,12,12,12,30,30,30,30,33,33,8,8,8,8,8,8},
						'{8,8,8,8,8,8,28,33,33,33,33,13,30,30,30,30,30,30,30,30,33,33,12,12,12,12,12,33,33,12,12,12,12,12,12,12,30,30,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,28,24,13,13,13,1,1,30,30,30,13,1,33,1,13,13,30,30,30,30,30,13,32,8,8,33,8,8,10,19,33,8,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,28,24,22,19,30,33,33,19,30,30,1,33,33,33,19,30,30,30,30,30,30,30,30,8,8,8,8,8,32,19,8,8,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,28,28,24,30,27,27,27,27,22,19,33,1,30,19,30,30,30,30,30,30,30,30,30,30,10,32,8,8,8,8,8,8,8,10,33,8,8,8,8,8,8},
						'{8,8,8,8,28,27,27,27,30,27,27,24,27,30,19,33,1,30,30,30,30,12,22,30,30,30,30,30,30,30,32,8,8,8,8,8,8,8,30,32,8,8,8,8,8,8},
						'{8,8,8,8,28,27,30,32,8,8,28,30,30,30,22,30,1,33,33,33,30,12,30,30,30,30,30,30,30,8,8,8,33,30,30,30,30,30,30,30,19,33,8,8,8,8},
						'{8,8,8,8,8,33,32,33,8,8,27,19,30,30,30,30,13,1,33,33,33,32,32,32,32,32,32,32,32,8,8,8,32,30,30,30,30,30,30,30,12,32,8,8,8,8},
						'{8,8,8,27,8,8,8,8,8,33,30,30,30,30,30,30,30,30,30,30,8,8,8,8,8,8,8,8,8,8,8,30,30,30,30,30,30,30,12,12,12,19,19,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,33,30,30,19,30,19,10,33,33,33,8,8,8,8,8,8,8,8,8,8,8,33,33,33,10,19,30,30,33,33,33,32,19,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,8,32,30,30,30,30,33,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,32,30,30,30,8,8,8,33,19,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8}};
		
		
		kraid_g = '{'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,33,25,8,8,8,8,25,33,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,21,33,8,8,8,21,32,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,8,8,8,21,32,8,8,8,32,21,8,8,21,32,31,31,31,31,31,8,8,31,8,8,8,31,8,8,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,8,8,8,32,32,8,8,8,32,21,8,8,21,25,30,30,30,30,32,8,8,8,8,8,33,32,8,8,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,21,33,8,32,21,31,32,15,21,21,21,21,21,21,15,32,33,16,21,21,15,8,8,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,8,8,33,33,32,33,8,8,31,21,30,30,21,21,21,3,16,21,21,21,21,31,35,21,10,33,33,33,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,8,25,21,21,30,33,28,13,25,21,21,21,21,21,21,31,33,3,21,21,21,21,21,21,33,33,35,21,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,25,31,32,32,30,30,27,33,33,30,21,21,21,21,21,35,33,28,13,33,33,33,16,21,21,21,35,35,33,8,25,33,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,15,21,0,13,13,13,13,33,16,21,21,21,21,21,21,10,33,28,13,33,33,33,33,21,21,21,21,21,33,33,21,32,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,15,30,13,33,33,33,33,21,21,21,33,33,33,33,21,21,21,16,33,25,21,21,30,33,16,21,21,21,21,21,21,32,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,33,10,30,27,33,33,33,33,21,21,3,16,33,33,33,35,35,21,31,33,10,30,30,25,33,16,25,21,21,21,21,25,33,8,8,8,8,8,8},
						'{8,8,8,31,8,8,15,32,13,28,33,33,33,33,33,21,31,33,3,21,21,21,33,16,21,21,21,33,33,13,28,33,33,33,3,21,21,21,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,32,30,13,28,28,33,16,16,33,33,33,16,35,21,10,31,16,3,21,21,21,31,16,28,28,33,33,28,3,21,21,21,8,8,8,8,8,8,8,8},
						'{8,8,8,8,31,31,31,31,13,13,13,30,21,21,32,8,33,21,21,21,33,33,21,21,21,21,21,21,21,33,33,33,33,13,25,21,21,25,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,8,33,30,30,30,30,33,8,33,21,21,21,33,33,16,33,16,33,16,35,21,3,3,3,25,25,21,21,21,21,32,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,8,33,15,32,31,31,31,8,33,21,21,21,33,33,33,33,33,33,33,32,21,21,21,21,21,21,21,21,21,21,21,32,8,8,8,8,8,8},
						'{8,8,8,8,25,25,15,33,8,8,8,31,31,8,8,8,8,8,32,21,35,3,33,33,33,16,25,8,8,21,21,21,21,21,21,21,21,21,21,32,8,8,8,8,8,8},
						'{8,8,8,8,32,30,21,32,8,8,8,8,31,8,8,8,8,8,33,21,21,21,33,33,33,3,15,8,8,25,21,21,21,21,21,21,21,21,21,32,8,8,8,8,8,8},
						'{8,8,32,15,32,13,13,32,21,33,8,8,8,8,8,8,8,8,8,8,25,21,21,21,21,21,21,8,8,8,8,21,21,21,21,21,21,21,21,21,15,33,8,8,8,8},
						'{8,8,33,30,13,13,13,30,30,8,8,8,8,8,8,8,8,8,8,8,33,32,32,32,32,32,32,33,8,8,8,32,25,21,21,21,3,3,21,21,21,33,8,8,8,8},
						'{8,8,8,13,13,13,13,13,13,13,13,31,13,8,8,21,33,8,8,8,8,8,8,8,8,8,8,32,21,8,8,8,33,21,21,21,33,33,21,21,21,33,8,8,8,8},
						'{8,33,33,13,13,13,13,31,8,8,8,8,8,8,8,21,25,33,33,33,32,33,33,33,8,8,8,33,33,33,33,8,33,21,21,21,3,31,21,21,21,33,8,8,8,8},
						'{33,15,30,13,13,13,13,8,8,8,8,8,8,8,8,15,21,21,21,21,21,21,21,32,8,8,8,8,8,21,32,8,33,15,21,21,15,21,21,21,21,33,8,8,8,8},
						'{28,30,13,13,33,33,25,33,8,8,8,8,8,25,25,21,21,21,21,21,21,21,21,21,32,32,32,32,25,8,8,8,8,8,8,8,21,21,21,32,8,8,8,8,8,8},
						'{33,13,13,13,33,33,21,32,8,8,8,8,8,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,8,8,8,8,8,8,8,25,21,21,32,8,8,8,8,8,8},
						'{33,33,28,13,25,21,21,32,31,31,31,8,8,8,8,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,15,8,8,8,8,8,8,8,8,8,8,8,8},
						'{33,33,28,13,21,21,30,30,13,13,31,8,8,8,8,21,21,21,21,21,21,21,21,21,35,3,35,21,21,21,21,21,21,15,33,8,8,8,8,8,8,8,8,8,8,8},
						'{33,33,33,33,25,30,13,13,13,13,31,8,8,21,21,21,21,21,21,21,21,21,21,10,33,33,33,3,21,21,21,21,21,21,21,15,21,21,8,8,8,8,8,8,8,8},
						'{33,33,33,16,30,30,13,13,13,31,8,8,8,33,32,21,21,21,21,21,3,31,3,33,33,33,16,35,21,21,21,21,21,21,21,15,32,33,8,8,8,8,8,8,8,8},
						'{33,33,3,21,13,13,13,13,31,8,8,8,8,8,8,21,21,21,21,21,33,33,33,33,33,16,21,21,21,21,21,21,21,21,21,15,8,8,8,8,8,8,8,8,8,8},
						'{33,3,30,30,13,13,13,31,8,8,8,33,32,8,8,21,21,21,21,21,10,3,33,33,33,33,16,33,16,21,21,21,21,21,31,33,32,33,8,8,8,8,8,8,8,8},
						'{16,21,30,31,31,13,31,8,8,8,8,32,21,8,8,21,21,21,21,21,21,21,33,33,33,33,33,33,33,21,21,21,21,21,33,33,35,25,8,8,8,8,8,8,8,8},
						'{8,31,13,31,8,8,8,8,8,33,25,33,8,25,32,8,33,21,21,21,21,21,35,35,35,35,25,33,33,33,33,33,33,33,31,21,21,21,25,33,8,8,8,8,8,8},
						'{8,31,31,31,8,8,8,8,8,33,25,8,33,21,25,8,33,21,25,21,21,21,21,21,21,21,21,33,33,33,33,33,33,33,3,21,21,21,21,32,8,8,8,8,8,8},
						'{8,8,8,13,25,25,31,8,8,8,8,32,21,21,25,8,8,8,8,8,8,8,21,3,33,33,33,3,21,21,35,33,33,33,3,21,21,21,21,21,15,33,8,8,8,8},
						'{8,8,33,30,10,25,13,8,8,8,8,33,32,32,33,8,8,8,8,8,8,8,32,33,33,33,33,35,21,3,31,16,33,33,16,3,3,3,3,35,21,33,8,8,8,8},
						'{8,8,32,21,13,13,13,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,21,30,13,25,21,33,33,21,10,33,33,33,33,33,33,33,21,33,8,8,8,8},
						'{8,8,8,30,13,13,28,8,8,8,8,33,33,33,33,33,33,33,33,33,8,8,33,32,30,27,28,33,16,31,10,10,31,33,33,16,16,16,33,33,21,33,8,8,8,8},
						'{8,8,8,31,31,13,33,33,13,8,8,32,21,21,21,21,21,21,21,21,8,8,15,30,13,28,33,33,33,21,30,13,28,33,3,21,21,21,33,8,15,33,8,8,8,8},
						'{8,8,8,8,31,13,30,25,25,32,25,21,21,33,33,33,33,33,3,21,25,32,8,33,33,33,33,31,35,30,27,33,31,3,21,21,21,21,3,32,8,8,8,8,8,8},
						'{8,8,8,8,31,13,0,21,21,21,21,21,21,33,33,33,33,33,3,21,21,21,33,33,33,33,33,35,30,13,13,33,16,21,21,21,21,21,21,32,8,8,8,8,8,8},
						'{8,8,8,31,8,33,21,30,13,13,13,13,13,33,33,21,16,33,33,33,35,21,21,21,21,21,21,33,33,33,33,21,21,21,21,21,21,21,21,21,21,33,8,8,8,8},
						'{8,8,8,31,8,33,30,30,13,13,13,27,13,33,16,21,3,33,33,33,21,21,21,21,35,35,3,33,33,33,33,21,21,21,21,21,21,21,21,21,25,33,8,8,8,8},
						'{8,8,8,8,31,13,13,13,13,28,33,33,33,21,21,21,21,21,21,21,21,21,21,3,33,33,33,33,33,33,33,21,21,21,21,21,21,21,21,32,8,8,8,8,8,8},
						'{8,8,8,8,8,8,13,13,28,33,33,33,16,21,21,21,21,21,21,21,3,31,21,35,16,16,16,33,33,16,10,21,21,21,21,21,21,21,33,33,8,8,8,8,8,8},
						'{8,8,8,8,8,8,31,28,33,33,33,3,21,21,21,21,21,21,21,21,33,33,21,21,21,21,21,33,33,21,21,21,21,21,21,21,21,21,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,31,13,3,3,3,16,16,21,21,21,3,16,33,16,3,3,21,21,21,21,21,3,32,8,8,33,8,8,25,15,33,8,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,31,30,21,21,21,33,33,21,21,21,31,33,33,33,35,21,21,21,21,21,21,21,21,8,8,8,8,8,32,15,8,8,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,31,31,30,21,25,13,13,13,21,35,33,16,21,25,21,21,21,21,21,21,21,21,21,21,25,32,8,8,8,8,8,8,8,25,33,8,8,8,8,8,8},
						'{8,8,8,8,31,13,13,32,15,32,13,13,13,21,35,33,31,21,30,21,30,21,21,21,21,21,21,21,21,21,32,8,8,8,8,8,8,8,21,32,8,8,8,8,8,8},
						'{8,8,8,8,31,13,21,32,8,8,31,30,21,21,21,21,31,33,33,33,21,21,21,21,21,21,21,21,21,8,8,8,33,21,21,21,21,21,21,21,15,33,8,8,8,8},
						'{8,8,8,8,8,33,32,33,8,8,32,21,21,21,21,21,3,16,33,33,33,32,32,32,32,32,32,32,32,8,8,8,32,21,21,21,21,21,21,21,21,32,8,8,8,8},
						'{8,8,8,13,8,8,8,8,8,33,21,21,21,21,21,21,21,21,21,21,8,8,8,8,8,8,8,8,8,8,8,21,21,21,21,21,21,21,21,21,21,15,15,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,33,21,21,21,21,21,25,33,33,33,8,8,8,8,8,8,8,8,8,8,8,33,33,33,25,21,21,21,33,33,33,32,15,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,8,32,21,21,21,21,33,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,32,21,21,21,8,8,8,33,15,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8},
						'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8}};
		
		
		kraid_n = '{'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,16,18,33,33,33,33,18,31,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,31,18,16,33,33,33,18,25,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,18,25,33,33,33,25,18,33,33,18,30,20,20,20,20,20,33,33,20,28,33,28,20,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,25,25,33,33,33,25,18,33,33,2,18,27,27,27,27,27,33,31,28,28,31,31,27,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,2,31,33,25,18,20,19,2,2,2,2,2,2,18,2,30,33,31,2,2,2,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,31,31,31,25,31,31,28,25,2,30,30,2,2,2,25,31,18,2,2,2,31,18,2,10,32,31,31,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,18,2,2,30,33,28,20,30,2,2,2,2,2,2,31,33,25,2,2,2,2,2,2,31,33,18,18,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,18,25,30,27,27,27,27,33,31,22,2,2,2,2,2,18,33,28,20,33,33,33,31,2,2,2,18,18,33,33,18,31,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,31,2,2,0,19,20,20,20,33,31,2,2,2,2,2,2,10,33,28,20,33,33,33,33,2,2,2,2,2,33,33,18,25,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,2,27,20,33,33,33,33,18,2,2,31,33,33,33,2,2,18,31,33,25,2,2,30,33,31,2,2,2,2,2,2,25,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,31,22,27,27,33,33,33,33,2,18,25,31,33,33,33,18,18,2,31,33,30,30,22,25,33,16,25,18,2,2,2,18,31,33,33,33,33,33,33},
						'{33,33,28,20,33,33,2,30,20,28,33,33,33,33,33,2,31,33,25,2,2,2,33,16,2,2,2,33,33,20,28,33,33,33,25,2,2,2,33,33,33,33,33,33,33,33},
						'{33,33,33,28,28,28,30,27,20,28,28,31,31,31,31,31,31,31,18,2,30,31,31,25,2,2,2,31,31,28,28,33,33,28,25,2,2,2,33,33,33,33,33,33,33,33},
						'{33,33,33,33,20,20,20,20,19,20,20,22,2,2,30,33,31,2,2,2,33,33,2,2,2,2,2,2,2,33,33,33,33,20,30,2,2,18,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,28,33,28,10,30,27,27,27,10,33,31,18,2,2,33,33,16,33,16,33,16,18,2,25,25,25,30,25,2,2,2,18,25,32,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,31,2,27,20,20,20,33,31,2,2,18,33,33,33,33,33,33,33,25,2,18,2,2,2,2,2,2,2,2,2,30,33,33,33,33,33,33},
						'{33,33,33,33,18,18,2,10,33,33,33,20,20,33,33,33,33,33,25,2,18,25,33,33,33,31,18,31,33,2,2,2,2,2,2,2,2,2,2,10,33,33,33,33,33,33},
						'{33,33,33,33,30,22,2,10,33,33,33,28,20,33,33,33,33,33,31,18,2,18,33,33,33,25,2,33,33,18,18,2,2,2,2,2,2,2,2,30,33,33,33,33,33,33},
						'{33,33,25,2,19,20,20,27,2,32,33,33,33,33,33,33,33,33,33,33,18,2,18,18,2,2,2,33,33,33,33,2,2,2,2,2,2,2,2,2,2,31,33,33,33,33},
						'{33,33,10,30,20,20,20,27,30,31,33,33,33,33,33,33,33,33,33,33,31,25,25,25,25,25,25,31,33,33,33,25,18,2,2,2,25,25,2,2,2,32,33,33,33,33},
						'{33,33,28,19,20,19,20,20,20,19,19,20,19,33,33,2,31,33,33,33,33,33,33,33,33,33,33,25,2,33,33,33,31,2,2,2,33,33,2,2,2,31,33,33,33,33},
						'{33,31,27,19,20,20,20,20,28,28,28,28,33,33,33,2,18,10,31,31,25,31,31,16,33,33,33,16,31,31,31,33,31,2,2,2,25,31,2,2,2,31,33,33,33,33},
						'{31,2,27,20,20,19,20,28,33,33,33,33,33,33,33,2,2,2,2,2,2,2,2,25,33,33,33,33,33,18,25,33,31,2,2,2,2,2,2,18,2,31,33,33,33,33},
						'{28,27,20,19,33,33,30,31,33,33,33,33,33,18,18,2,2,2,2,2,2,2,2,18,25,25,25,25,18,33,33,33,33,33,33,33,18,2,2,25,33,33,33,33,33,33},
						'{33,19,20,20,33,33,2,25,33,33,33,33,33,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,33,33,33,33,33,33,33,18,2,2,25,33,33,33,33,33,33},
						'{33,33,28,19,18,2,2,30,20,20,20,33,33,33,33,2,2,2,2,2,2,2,2,2,2,2,2,2,18,18,18,18,2,2,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,28,20,2,2,22,30,20,20,20,33,33,33,31,2,2,2,2,2,2,2,2,18,18,25,18,18,2,2,2,2,2,2,32,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,18,22,20,20,20,19,20,33,33,18,2,2,2,2,2,2,2,2,2,30,33,33,33,25,2,2,2,2,2,2,2,2,2,18,33,33,33,33,33,33,33,33},
						'{33,33,33,31,30,30,20,20,20,20,28,33,33,31,25,2,2,2,2,2,25,31,25,31,33,33,31,18,2,2,2,2,2,2,2,2,25,31,33,33,33,33,33,33,33,33},
						'{33,33,25,2,20,20,20,19,20,28,33,33,33,33,33,2,18,2,2,2,33,33,33,33,33,31,2,2,2,2,2,2,2,2,2,2,33,33,33,33,33,33,33,33,33,33},
						'{33,25,27,27,19,20,20,20,33,33,33,31,25,33,33,2,2,2,2,2,10,25,33,33,33,33,16,31,16,2,2,2,18,2,31,16,25,31,33,33,33,33,33,33,33,33},
						'{31,2,27,20,20,19,20,28,33,33,33,25,18,33,33,2,2,2,2,2,2,2,33,33,33,33,33,33,33,18,2,2,2,2,31,33,18,18,33,33,33,33,33,33,33,33},
						'{28,20,19,20,33,33,33,33,33,31,18,16,33,18,25,33,31,2,2,2,2,2,18,18,18,18,18,33,33,33,33,33,33,33,31,18,18,2,18,31,33,33,33,33,33,33},
						'{33,20,20,20,33,33,33,33,33,31,18,33,33,2,18,33,16,18,18,18,18,18,2,18,18,2,2,33,33,33,33,33,33,33,25,18,2,2,2,25,33,33,33,33,33,33},
						'{33,33,28,19,18,18,20,28,33,33,33,25,2,18,18,33,33,33,33,33,33,33,2,25,33,33,33,25,2,18,18,33,33,33,25,2,2,2,2,2,2,31,33,33,33,33},
						'{33,33,1,27,10,30,20,28,33,33,33,31,25,25,31,33,33,33,33,33,33,33,25,31,31,33,33,18,2,25,31,16,33,33,16,25,25,25,25,18,2,32,33,33,33,33},
						'{33,33,25,18,19,20,20,28,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,31,2,27,19,30,2,33,33,2,10,33,33,33,33,33,33,33,2,32,33,33,33,33},
						'{33,33,31,27,20,20,28,28,28,33,33,16,31,31,31,31,31,31,31,31,33,33,31,10,27,27,28,31,31,31,10,10,1,33,33,31,31,31,33,31,2,32,33,33,33,33},
						'{33,33,28,20,20,20,33,33,19,28,33,25,2,2,2,2,2,2,2,2,33,33,2,30,20,28,33,33,33,2,22,20,28,33,25,2,2,18,33,33,2,32,33,33,33,33},
						'{33,33,33,33,20,20,30,18,30,30,18,2,2,33,33,33,33,33,25,2,18,25,33,33,33,33,33,31,18,27,27,33,31,25,18,2,2,18,25,25,33,33,33,33,33,33},
						'{33,33,33,33,20,19,0,2,2,2,2,2,2,33,33,33,33,33,25,2,18,18,33,33,33,33,33,18,22,19,20,33,31,2,2,2,2,2,2,25,33,33,33,33,33,33},
						'{33,33,28,20,33,33,2,30,20,20,20,20,20,33,33,18,31,33,33,33,18,2,18,18,18,18,2,33,33,33,33,18,2,2,2,18,2,2,2,18,18,31,33,33,33,33},
						'{33,33,28,20,33,33,22,30,20,20,20,27,20,33,16,2,25,33,33,33,18,2,2,18,18,18,25,33,33,33,33,2,2,2,2,2,2,18,2,18,18,16,33,33,33,33},
						'{33,33,33,33,20,20,20,20,20,28,33,33,33,2,2,2,2,2,2,2,2,2,2,25,33,33,33,33,33,33,33,2,2,2,2,2,2,2,2,25,33,33,33,33,33,33},
						'{33,33,33,33,28,28,19,20,28,33,33,33,31,2,2,2,2,2,2,2,25,31,2,18,31,31,31,33,33,31,10,2,2,2,2,2,2,18,31,16,33,33,33,33,33,33},
						'{33,33,33,33,33,33,20,28,33,33,33,25,2,2,2,2,2,2,2,2,33,33,2,2,2,2,2,33,33,2,2,2,2,2,2,2,2,18,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,20,19,25,25,25,31,16,2,2,2,25,16,31,16,25,25,2,2,2,2,2,25,25,31,31,32,31,31,18,2,31,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,20,27,2,18,2,33,33,18,2,2,31,33,33,33,18,2,2,2,2,2,2,2,2,33,33,33,33,33,30,2,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,28,20,20,27,2,25,20,20,20,2,18,33,31,2,18,2,2,2,2,2,2,2,2,2,2,18,25,33,33,33,33,33,33,33,18,31,33,33,33,33,33,33},
						'{33,33,33,33,20,20,20,27,2,27,20,19,20,2,18,33,31,2,30,2,22,2,2,2,2,2,2,2,18,18,25,33,33,33,33,33,33,33,2,25,33,33,33,33,33,33},
						'{33,33,33,33,20,20,2,25,33,28,20,30,2,2,2,2,31,33,33,33,2,2,2,2,2,2,2,2,2,33,33,33,16,18,2,18,18,2,2,2,2,31,33,33,33,33},
						'{33,33,33,33,28,27,25,31,33,33,27,18,2,2,2,2,25,16,33,16,10,30,25,25,25,25,25,25,25,33,33,33,25,2,2,2,2,2,2,2,2,30,33,33,33,33},
						'{33,33,28,19,33,33,33,33,33,31,2,2,2,2,2,2,2,2,2,2,33,33,33,33,33,33,33,33,33,33,33,2,2,2,2,2,2,2,2,2,2,2,2,33,33,33},
						'{33,33,33,28,33,33,33,33,33,33,31,18,2,18,2,18,18,31,31,31,33,33,33,33,33,33,33,33,33,33,33,31,31,31,18,18,2,18,32,32,32,30,2,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,25,2,2,2,2,31,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,25,2,2,18,33,33,33,31,2,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33}};
						
						shoot =   '{'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
										'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
										'{33,33,33,33,31,31,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
										'{33,33,33,33,18,18,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
										'{33,33,33,33,18,2,25,31,33,33,33,33,33,33,33,25,31,33,33,33,33},
										'{33,33,33,33,18,2,2,25,33,33,33,33,33,33,33,2,31,33,33,33,33},
										'{33,33,33,33,2,2,2,2,2,16,33,33,33,18,2,2,2,2,33,33,33},
										'{33,33,33,33,30,30,2,2,2,31,33,33,33,2,2,2,2,2,33,33,33},
										'{33,33,33,33,33,33,2,2,2,2,2,2,2,2,2,2,2,2,33,33,33},
										'{33,33,33,33,33,33,2,2,2,2,2,2,2,2,2,2,2,2,33,33,33},
										'{33,33,33,33,33,33,0,2,2,2,2,2,2,2,2,2,2,2,32,33,33},
										'{33,33,33,33,33,33,31,25,2,2,2,2,2,2,2,2,10,32,33,33,33},
										'{33,33,33,33,33,33,33,33,2,2,2,2,2,2,2,2,25,33,33,33,33},
										'{33,33,33,33,33,33,33,33,33,33,33,2,2,2,30,33,33,33,33,33,33},
										'{33,33,33,33,33,33,33,33,33,33,33,10,2,2,30,33,33,33,33,33,33},
										'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
										'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
										'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33}};
										
						attack =  '{'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
										'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
										'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
										'{33,33,33,31,33,31,33,31,33,31,33,33,33,33,33,33,33},
										'{33,33,2,2,2,2,2,2,2,2,2,33,33,33,33,33,33},
										'{33,33,32,32,32,32,32,32,32,32,32,28,28,28,28,28,33},
										'{33,33,33,33,33,33,33,33,33,33,33,20,20,20,20,20,33},
										'{33,33,25,25,25,25,25,25,25,25,25,33,33,33,33,33,33},
										'{33,33,18,2,2,2,2,2,2,2,18,33,33,33,33,33,33},
										'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
										'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
										'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33}};
	end
	
	always_comb begin
		// Defaults:
		draw = 0;
		color = 0;

		if(vga_x >= kraid_x && vga_x < kraid_x + kraid_w && vga_y >= kraid_y && vga_y < kraid_y + kraid_h && kraid_g_en) begin
			if(kraid_g[vga_y - kraid_y][vga_x - kraid_x] != 8) begin
				draw = 1'b1;
				color = kraid_g[vga_y - kraid_y][vga_x - kraid_x];
			end
			if(kraid_dir == 1'b1) begin
				if(kraid_g[vga_y - kraid_y][kraid_x + kraid_w - 1 - vga_x] != 8) begin
					draw = 1'b1;
					color = kraid_g[vga_y - kraid_y][kraid_x + kraid_w - 1 - vga_x];
				end
			end
		end
		if(vga_x >= kraid_x && vga_x < kraid_x + kraid_w && vga_y >= kraid_y && vga_y < kraid_y + kraid_h && kraid_r_en) begin
			if(kraid_r[vga_y - kraid_y][vga_x - kraid_x] != 8) begin
				draw = 1'b1;
				color = kraid_r[vga_y - kraid_y][vga_x - kraid_x];
			end
			if(kraid_dir == 1'b1) begin
				if(kraid_r[vga_y - kraid_y][kraid_x + kraid_w - 1 - vga_x] != 8) begin
					draw = 1'b1;
					color = kraid_r[vga_y - kraid_y][kraid_x + kraid_w - 1 - vga_x];
				end
			end
		end
		if(vga_x >= kraid_x && vga_x < kraid_x + kraid_w && vga_y >= kraid_y && vga_y < kraid_y + kraid_h && kraid_n_en) begin
			if(kraid_n[vga_y - kraid_y][vga_x - kraid_x] != 33) begin
				draw = 1'b1;
				color = kraid_n[vga_y - kraid_y][vga_x - kraid_x];
			end
			if(kraid_dir == 1'b1) begin
				if(kraid_n[vga_y - kraid_y][kraid_x + kraid_w - 1 - vga_x] != 33) begin
					draw = 1'b1;
					color = kraid_n[vga_y - kraid_y][kraid_x + kraid_w - 1 - vga_x];
				end
			end
		end
		// Shoot:
		if(vga_x >= shoot_x && vga_x < shoot_x + shoot_w && vga_y >= shoot_y && vga_y < shoot_y + shoot_h && kraid_shoot_en) begin
			if(shoot[vga_y - shoot_y][vga_x - shoot_x] != 33) begin
				draw = 1'b1;
				color = shoot[vga_y - shoot_y][vga_x - shoot_x];
			end
			if(kraid_as_dir == 1'b1) begin
				if(shoot[vga_y - shoot_y][shoot_x + shoot_w - 1 - vga_x] != 33) begin
					draw = 1'b1;
					color = shoot[vga_y - shoot_y][shoot_x + shoot_w - 1 - vga_x];
				end
			end
		end
		// Throw:
		if(vga_x >= throw_x && vga_x < throw_x + attack_w && vga_y >= throw_y && vga_y < throw_y + attack_h && kraid_throw_en) begin
			if(attack[vga_y - throw_y][vga_x - throw_x] != 33) begin
				draw = 1'b1;
				color = attack[vga_y - throw_y][vga_x - throw_x];
			end
			if(kraid_as_dir == 1'b1) begin
				if(attack[vga_y - throw_y][throw_x + attack_w - 1 - vga_x] != 33) begin
					draw = 1'b1;
					color = attack[vga_y - throw_y][throw_x + attack_w - 1 - vga_x];
				end
			end
		end
		// Throw2:
		if(vga_x >= throw_2_x && vga_x < throw_2_x + attack_w && vga_y >= throw_2_y && vga_y < throw_2_y + attack_h && kraid_throw_2_en) begin
			if(attack[vga_y - throw_2_y][vga_x - throw_2_x] != 33) begin
				draw = 1'b1;
				color = attack[vga_y - throw_2_y][vga_x - throw_2_x];
			end
			if(kraid_as_dir == 1'b1) begin
				if(attack[vga_y - throw_2_y][throw_2_x + attack_w - 1 - vga_x] != 33) begin
					draw = 1'b1;
					color = attack[vga_y - throw_2_y][throw_2_x + attack_w - 1 - vga_x];
				end
			end
		end
	end
endmodule