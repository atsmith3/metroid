// nios_system.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module nios_system (
		output wire        bullet1_en_export,      //      bullet1_en.export
		output wire [9:0]  bullet1_x_export,       //       bullet1_x.export
		output wire [9:0]  bullet1_y_export,       //       bullet1_y.export
		output wire        bullet2_en_export,      //      bullet2_en.export
		output wire [9:0]  bullet2_x_export,       //       bullet2_x.export
		output wire [9:0]  bullet2_y_export,       //       bullet2_y.export
		output wire        bullet3_en_export,      //      bullet3_en.export
		output wire [9:0]  bullet3_x_export,       //       bullet3_x.export
		output wire [9:0]  bullet3_y_export,       //       bullet3_y.export
		input  wire        clk_clk,                //             clk.clk
		output wire        explosion1_en_export,   //   explosion1_en.export
		output wire [9:0]  explosion1_x_export,    //    explosion1_x.export
		output wire [9:0]  explosion1_y_export,    //    explosion1_y.export
		output wire        explosion2_en_export,   //   explosion2_en.export
		output wire [9:0]  explosion2_x_export,    //    explosion2_x.export
		output wire [9:0]  explosion2_y_export,    //    explosion2_y.export
		output wire        explosion3_en_export,   //   explosion3_en.export
		output wire [9:0]  explosion3_x_export,    //    explosion3_x.export
		output wire [9:0]  explosion3_y_export,    //    explosion3_y.export
		output wire [1:0]  health_export,          //          health.export
		input  wire [1:0]  key_export,             //             key.export
		output wire [15:0] keycode_export,         //         keycode.export
		output wire        loss_en_export,         //         loss_en.export
		output wire        monster1_en_export,     //     monster1_en.export
		output wire [9:0]  monster1_x_export,      //      monster1_x.export
		output wire [9:0]  monster1_y_export,      //      monster1_y.export
		output wire        monster2_en_export,     //     monster2_en.export
		output wire [9:0]  monster2_x_export,      //      monster2_x.export
		output wire [9:0]  monster2_y_export,      //      monster2_y.export
		output wire        monster3_en_export,     //     monster3_en.export
		output wire [9:0]  monster3_x_export,      //      monster3_x.export
		output wire [9:0]  monster3_y_export,      //      monster3_y.export
		output wire [1:0]  otg_hpi_address_export, // otg_hpi_address.export
		output wire        otg_hpi_cs_export,      //      otg_hpi_cs.export
		input  wire [15:0] otg_hpi_data_in_port,   //    otg_hpi_data.in_port
		output wire [15:0] otg_hpi_data_out_port,  //                .out_port
		output wire        otg_hpi_r_export,       //       otg_hpi_r.export
		output wire        otg_hpi_w_export,       //       otg_hpi_w.export
		input  wire        reset_reset_n,          //           reset.reset_n
		output wire        samus_dir_export,       //       samus_dir.export
		output wire        samus_en_export,        //        samus_en.export
		output wire        samus_jump_export,      //      samus_jump.export
		output wire        samus_walk_export,      //      samus_walk.export
		output wire [9:0]  samus_x_export,         //         samus_x.export
		output wire [9:0]  samus_y_export,         //         samus_y.export
		output wire [2:0]  scene_sel_export,       //       scene_sel.export
		output wire        sdram_clk_clk,          //       sdram_clk.clk
		output wire [12:0] sdram_wire_addr,        //      sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,          //                .ba
		output wire        sdram_wire_cas_n,       //                .cas_n
		output wire        sdram_wire_cke,         //                .cke
		output wire        sdram_wire_cs_n,        //                .cs_n
		inout  wire [31:0] sdram_wire_dq,          //                .dq
		output wire [3:0]  sdram_wire_dqm,         //                .dqm
		output wire        sdram_wire_ras_n,       //                .ras_n
		output wire        sdram_wire_we_n,        //                .we_n
		output wire        title_en_export,        //        title_en.export
		output wire        win_en_export           //          win_en.export
	);

	wire         sdram_pll_c0_clk;                                            // sdram_pll:c0 -> [mm_interconnect_0:sdram_pll_c0_clk, rst_controller_001:clk, sdram:clk]
	wire  [31:0] nios2_qsys_0_data_master_readdata;                           // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire         nios2_qsys_0_data_master_debugaccess;                        // nios2_qsys_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire  [28:0] nios2_qsys_0_data_master_address;                            // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                         // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire         nios2_qsys_0_data_master_read;                               // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire         nios2_qsys_0_data_master_write;                              // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire  [31:0] nios2_qsys_0_data_master_writedata;                          // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         nios2_qsys_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [28:0] nios2_qsys_0_instruction_master_address;                     // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                        // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;       // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;        // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_readdata;     // nios2_qsys_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_qsys_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_waitrequest;  // nios2_qsys_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_qsys_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_debugaccess -> nios2_qsys_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_address -> nios2_qsys_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_read -> nios2_qsys_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_byteenable -> nios2_qsys_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_write -> nios2_qsys_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_writedata -> nios2_qsys_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_readdata;              // sdram_pll:readdata -> mm_interconnect_0:sdram_pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_sdram_pll_pll_slave_address;               // mm_interconnect_0:sdram_pll_pll_slave_address -> sdram_pll:address
	wire         mm_interconnect_0_sdram_pll_pll_slave_read;                  // mm_interconnect_0:sdram_pll_pll_slave_read -> sdram_pll:read
	wire         mm_interconnect_0_sdram_pll_pll_slave_write;                 // mm_interconnect_0:sdram_pll_pll_slave_write -> sdram_pll:write
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_writedata;             // mm_interconnect_0:sdram_pll_pll_slave_writedata -> sdram_pll:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [1:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_otg_hpi_address_s1_chipselect;             // mm_interconnect_0:otg_hpi_address_s1_chipselect -> otg_hpi_address:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_address_s1_readdata;               // otg_hpi_address:readdata -> mm_interconnect_0:otg_hpi_address_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_address_s1_address;                // mm_interconnect_0:otg_hpi_address_s1_address -> otg_hpi_address:address
	wire         mm_interconnect_0_otg_hpi_address_s1_write;                  // mm_interconnect_0:otg_hpi_address_s1_write -> otg_hpi_address:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_address_s1_writedata;              // mm_interconnect_0:otg_hpi_address_s1_writedata -> otg_hpi_address:writedata
	wire         mm_interconnect_0_otg_hpi_data_s1_chipselect;                // mm_interconnect_0:otg_hpi_data_s1_chipselect -> otg_hpi_data:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_data_s1_readdata;                  // otg_hpi_data:readdata -> mm_interconnect_0:otg_hpi_data_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_data_s1_address;                   // mm_interconnect_0:otg_hpi_data_s1_address -> otg_hpi_data:address
	wire         mm_interconnect_0_otg_hpi_data_s1_write;                     // mm_interconnect_0:otg_hpi_data_s1_write -> otg_hpi_data:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_data_s1_writedata;                 // mm_interconnect_0:otg_hpi_data_s1_writedata -> otg_hpi_data:writedata
	wire         mm_interconnect_0_otg_hpi_r_s1_chipselect;                   // mm_interconnect_0:otg_hpi_r_s1_chipselect -> otg_hpi_r:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_r_s1_readdata;                     // otg_hpi_r:readdata -> mm_interconnect_0:otg_hpi_r_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_r_s1_address;                      // mm_interconnect_0:otg_hpi_r_s1_address -> otg_hpi_r:address
	wire         mm_interconnect_0_otg_hpi_r_s1_write;                        // mm_interconnect_0:otg_hpi_r_s1_write -> otg_hpi_r:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_r_s1_writedata;                    // mm_interconnect_0:otg_hpi_r_s1_writedata -> otg_hpi_r:writedata
	wire         mm_interconnect_0_otg_hpi_w_s1_chipselect;                   // mm_interconnect_0:otg_hpi_w_s1_chipselect -> otg_hpi_w:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_w_s1_readdata;                     // otg_hpi_w:readdata -> mm_interconnect_0:otg_hpi_w_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_w_s1_address;                      // mm_interconnect_0:otg_hpi_w_s1_address -> otg_hpi_w:address
	wire         mm_interconnect_0_otg_hpi_w_s1_write;                        // mm_interconnect_0:otg_hpi_w_s1_write -> otg_hpi_w:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_w_s1_writedata;                    // mm_interconnect_0:otg_hpi_w_s1_writedata -> otg_hpi_w:writedata
	wire         mm_interconnect_0_otg_hpi_cs_s1_chipselect;                  // mm_interconnect_0:otg_hpi_cs_s1_chipselect -> otg_hpi_cs:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_cs_s1_readdata;                    // otg_hpi_cs:readdata -> mm_interconnect_0:otg_hpi_cs_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_cs_s1_address;                     // mm_interconnect_0:otg_hpi_cs_s1_address -> otg_hpi_cs:address
	wire         mm_interconnect_0_otg_hpi_cs_s1_write;                       // mm_interconnect_0:otg_hpi_cs_s1_write -> otg_hpi_cs:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_cs_s1_writedata;                   // mm_interconnect_0:otg_hpi_cs_s1_writedata -> otg_hpi_cs:writedata
	wire         mm_interconnect_0_keycode_s1_chipselect;                     // mm_interconnect_0:keycode_s1_chipselect -> keycode:chipselect
	wire  [31:0] mm_interconnect_0_keycode_s1_readdata;                       // keycode:readdata -> mm_interconnect_0:keycode_s1_readdata
	wire   [1:0] mm_interconnect_0_keycode_s1_address;                        // mm_interconnect_0:keycode_s1_address -> keycode:address
	wire         mm_interconnect_0_keycode_s1_write;                          // mm_interconnect_0:keycode_s1_write -> keycode:write_n
	wire  [31:0] mm_interconnect_0_keycode_s1_writedata;                      // mm_interconnect_0:keycode_s1_writedata -> keycode:writedata
	wire         mm_interconnect_0_key_s1_chipselect;                         // mm_interconnect_0:key_s1_chipselect -> key:chipselect
	wire  [31:0] mm_interconnect_0_key_s1_readdata;                           // key:readdata -> mm_interconnect_0:key_s1_readdata
	wire   [1:0] mm_interconnect_0_key_s1_address;                            // mm_interconnect_0:key_s1_address -> key:address
	wire         mm_interconnect_0_key_s1_write;                              // mm_interconnect_0:key_s1_write -> key:write_n
	wire  [31:0] mm_interconnect_0_key_s1_writedata;                          // mm_interconnect_0:key_s1_writedata -> key:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                       // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                         // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                      // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                          // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                             // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                       // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                    // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                            // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                        // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_samus_en_s1_chipselect;                    // mm_interconnect_0:samus_en_s1_chipselect -> samus_en:chipselect
	wire  [31:0] mm_interconnect_0_samus_en_s1_readdata;                      // samus_en:readdata -> mm_interconnect_0:samus_en_s1_readdata
	wire   [1:0] mm_interconnect_0_samus_en_s1_address;                       // mm_interconnect_0:samus_en_s1_address -> samus_en:address
	wire         mm_interconnect_0_samus_en_s1_write;                         // mm_interconnect_0:samus_en_s1_write -> samus_en:write_n
	wire  [31:0] mm_interconnect_0_samus_en_s1_writedata;                     // mm_interconnect_0:samus_en_s1_writedata -> samus_en:writedata
	wire         mm_interconnect_0_samus_x_s1_chipselect;                     // mm_interconnect_0:samus_x_s1_chipselect -> samus_x:chipselect
	wire  [31:0] mm_interconnect_0_samus_x_s1_readdata;                       // samus_x:readdata -> mm_interconnect_0:samus_x_s1_readdata
	wire   [1:0] mm_interconnect_0_samus_x_s1_address;                        // mm_interconnect_0:samus_x_s1_address -> samus_x:address
	wire         mm_interconnect_0_samus_x_s1_write;                          // mm_interconnect_0:samus_x_s1_write -> samus_x:write_n
	wire  [31:0] mm_interconnect_0_samus_x_s1_writedata;                      // mm_interconnect_0:samus_x_s1_writedata -> samus_x:writedata
	wire         mm_interconnect_0_samus_y_s1_chipselect;                     // mm_interconnect_0:samus_y_s1_chipselect -> samus_y:chipselect
	wire  [31:0] mm_interconnect_0_samus_y_s1_readdata;                       // samus_y:readdata -> mm_interconnect_0:samus_y_s1_readdata
	wire   [1:0] mm_interconnect_0_samus_y_s1_address;                        // mm_interconnect_0:samus_y_s1_address -> samus_y:address
	wire         mm_interconnect_0_samus_y_s1_write;                          // mm_interconnect_0:samus_y_s1_write -> samus_y:write_n
	wire  [31:0] mm_interconnect_0_samus_y_s1_writedata;                      // mm_interconnect_0:samus_y_s1_writedata -> samus_y:writedata
	wire         mm_interconnect_0_samus_walk_s1_chipselect;                  // mm_interconnect_0:samus_walk_s1_chipselect -> samus_walk:chipselect
	wire  [31:0] mm_interconnect_0_samus_walk_s1_readdata;                    // samus_walk:readdata -> mm_interconnect_0:samus_walk_s1_readdata
	wire   [1:0] mm_interconnect_0_samus_walk_s1_address;                     // mm_interconnect_0:samus_walk_s1_address -> samus_walk:address
	wire         mm_interconnect_0_samus_walk_s1_write;                       // mm_interconnect_0:samus_walk_s1_write -> samus_walk:write_n
	wire  [31:0] mm_interconnect_0_samus_walk_s1_writedata;                   // mm_interconnect_0:samus_walk_s1_writedata -> samus_walk:writedata
	wire         mm_interconnect_0_samus_jump_s1_chipselect;                  // mm_interconnect_0:samus_jump_s1_chipselect -> samus_jump:chipselect
	wire  [31:0] mm_interconnect_0_samus_jump_s1_readdata;                    // samus_jump:readdata -> mm_interconnect_0:samus_jump_s1_readdata
	wire   [1:0] mm_interconnect_0_samus_jump_s1_address;                     // mm_interconnect_0:samus_jump_s1_address -> samus_jump:address
	wire         mm_interconnect_0_samus_jump_s1_write;                       // mm_interconnect_0:samus_jump_s1_write -> samus_jump:write_n
	wire  [31:0] mm_interconnect_0_samus_jump_s1_writedata;                   // mm_interconnect_0:samus_jump_s1_writedata -> samus_jump:writedata
	wire         mm_interconnect_0_monster1_en_s1_chipselect;                 // mm_interconnect_0:monster1_en_s1_chipselect -> monster1_en:chipselect
	wire  [31:0] mm_interconnect_0_monster1_en_s1_readdata;                   // monster1_en:readdata -> mm_interconnect_0:monster1_en_s1_readdata
	wire   [1:0] mm_interconnect_0_monster1_en_s1_address;                    // mm_interconnect_0:monster1_en_s1_address -> monster1_en:address
	wire         mm_interconnect_0_monster1_en_s1_write;                      // mm_interconnect_0:monster1_en_s1_write -> monster1_en:write_n
	wire  [31:0] mm_interconnect_0_monster1_en_s1_writedata;                  // mm_interconnect_0:monster1_en_s1_writedata -> monster1_en:writedata
	wire         mm_interconnect_0_monster1_x_s1_chipselect;                  // mm_interconnect_0:monster1_x_s1_chipselect -> monster1_x:chipselect
	wire  [31:0] mm_interconnect_0_monster1_x_s1_readdata;                    // monster1_x:readdata -> mm_interconnect_0:monster1_x_s1_readdata
	wire   [1:0] mm_interconnect_0_monster1_x_s1_address;                     // mm_interconnect_0:monster1_x_s1_address -> monster1_x:address
	wire         mm_interconnect_0_monster1_x_s1_write;                       // mm_interconnect_0:monster1_x_s1_write -> monster1_x:write_n
	wire  [31:0] mm_interconnect_0_monster1_x_s1_writedata;                   // mm_interconnect_0:monster1_x_s1_writedata -> monster1_x:writedata
	wire         mm_interconnect_0_monster1_y_s1_chipselect;                  // mm_interconnect_0:monster1_y_s1_chipselect -> monster1_y:chipselect
	wire  [31:0] mm_interconnect_0_monster1_y_s1_readdata;                    // monster1_y:readdata -> mm_interconnect_0:monster1_y_s1_readdata
	wire   [1:0] mm_interconnect_0_monster1_y_s1_address;                     // mm_interconnect_0:monster1_y_s1_address -> monster1_y:address
	wire         mm_interconnect_0_monster1_y_s1_write;                       // mm_interconnect_0:monster1_y_s1_write -> monster1_y:write_n
	wire  [31:0] mm_interconnect_0_monster1_y_s1_writedata;                   // mm_interconnect_0:monster1_y_s1_writedata -> monster1_y:writedata
	wire         mm_interconnect_0_monster2_en_s1_chipselect;                 // mm_interconnect_0:monster2_en_s1_chipselect -> monster2_en:chipselect
	wire  [31:0] mm_interconnect_0_monster2_en_s1_readdata;                   // monster2_en:readdata -> mm_interconnect_0:monster2_en_s1_readdata
	wire   [1:0] mm_interconnect_0_monster2_en_s1_address;                    // mm_interconnect_0:monster2_en_s1_address -> monster2_en:address
	wire         mm_interconnect_0_monster2_en_s1_write;                      // mm_interconnect_0:monster2_en_s1_write -> monster2_en:write_n
	wire  [31:0] mm_interconnect_0_monster2_en_s1_writedata;                  // mm_interconnect_0:monster2_en_s1_writedata -> monster2_en:writedata
	wire         mm_interconnect_0_monster2_x_s1_chipselect;                  // mm_interconnect_0:monster2_x_s1_chipselect -> monster2_x:chipselect
	wire  [31:0] mm_interconnect_0_monster2_x_s1_readdata;                    // monster2_x:readdata -> mm_interconnect_0:monster2_x_s1_readdata
	wire   [1:0] mm_interconnect_0_monster2_x_s1_address;                     // mm_interconnect_0:monster2_x_s1_address -> monster2_x:address
	wire         mm_interconnect_0_monster2_x_s1_write;                       // mm_interconnect_0:monster2_x_s1_write -> monster2_x:write_n
	wire  [31:0] mm_interconnect_0_monster2_x_s1_writedata;                   // mm_interconnect_0:monster2_x_s1_writedata -> monster2_x:writedata
	wire         mm_interconnect_0_monster2_y_s1_chipselect;                  // mm_interconnect_0:monster2_y_s1_chipselect -> monster2_y:chipselect
	wire  [31:0] mm_interconnect_0_monster2_y_s1_readdata;                    // monster2_y:readdata -> mm_interconnect_0:monster2_y_s1_readdata
	wire   [1:0] mm_interconnect_0_monster2_y_s1_address;                     // mm_interconnect_0:monster2_y_s1_address -> monster2_y:address
	wire         mm_interconnect_0_monster2_y_s1_write;                       // mm_interconnect_0:monster2_y_s1_write -> monster2_y:write_n
	wire  [31:0] mm_interconnect_0_monster2_y_s1_writedata;                   // mm_interconnect_0:monster2_y_s1_writedata -> monster2_y:writedata
	wire         mm_interconnect_0_monster3_en_s1_chipselect;                 // mm_interconnect_0:monster3_en_s1_chipselect -> monster3_en:chipselect
	wire  [31:0] mm_interconnect_0_monster3_en_s1_readdata;                   // monster3_en:readdata -> mm_interconnect_0:monster3_en_s1_readdata
	wire   [1:0] mm_interconnect_0_monster3_en_s1_address;                    // mm_interconnect_0:monster3_en_s1_address -> monster3_en:address
	wire         mm_interconnect_0_monster3_en_s1_write;                      // mm_interconnect_0:monster3_en_s1_write -> monster3_en:write_n
	wire  [31:0] mm_interconnect_0_monster3_en_s1_writedata;                  // mm_interconnect_0:monster3_en_s1_writedata -> monster3_en:writedata
	wire         mm_interconnect_0_monster3_x_s1_chipselect;                  // mm_interconnect_0:monster3_x_s1_chipselect -> monster3_x:chipselect
	wire  [31:0] mm_interconnect_0_monster3_x_s1_readdata;                    // monster3_x:readdata -> mm_interconnect_0:monster3_x_s1_readdata
	wire   [1:0] mm_interconnect_0_monster3_x_s1_address;                     // mm_interconnect_0:monster3_x_s1_address -> monster3_x:address
	wire         mm_interconnect_0_monster3_x_s1_write;                       // mm_interconnect_0:monster3_x_s1_write -> monster3_x:write_n
	wire  [31:0] mm_interconnect_0_monster3_x_s1_writedata;                   // mm_interconnect_0:monster3_x_s1_writedata -> monster3_x:writedata
	wire         mm_interconnect_0_monster3_y_s1_chipselect;                  // mm_interconnect_0:monster3_y_s1_chipselect -> monster3_y:chipselect
	wire  [31:0] mm_interconnect_0_monster3_y_s1_readdata;                    // monster3_y:readdata -> mm_interconnect_0:monster3_y_s1_readdata
	wire   [1:0] mm_interconnect_0_monster3_y_s1_address;                     // mm_interconnect_0:monster3_y_s1_address -> monster3_y:address
	wire         mm_interconnect_0_monster3_y_s1_write;                       // mm_interconnect_0:monster3_y_s1_write -> monster3_y:write_n
	wire  [31:0] mm_interconnect_0_monster3_y_s1_writedata;                   // mm_interconnect_0:monster3_y_s1_writedata -> monster3_y:writedata
	wire         mm_interconnect_0_explosion1_en_s1_chipselect;               // mm_interconnect_0:explosion1_en_s1_chipselect -> explosion1_en:chipselect
	wire  [31:0] mm_interconnect_0_explosion1_en_s1_readdata;                 // explosion1_en:readdata -> mm_interconnect_0:explosion1_en_s1_readdata
	wire   [1:0] mm_interconnect_0_explosion1_en_s1_address;                  // mm_interconnect_0:explosion1_en_s1_address -> explosion1_en:address
	wire         mm_interconnect_0_explosion1_en_s1_write;                    // mm_interconnect_0:explosion1_en_s1_write -> explosion1_en:write_n
	wire  [31:0] mm_interconnect_0_explosion1_en_s1_writedata;                // mm_interconnect_0:explosion1_en_s1_writedata -> explosion1_en:writedata
	wire         mm_interconnect_0_explosion1_x_s1_chipselect;                // mm_interconnect_0:explosion1_x_s1_chipselect -> explosion1_x:chipselect
	wire  [31:0] mm_interconnect_0_explosion1_x_s1_readdata;                  // explosion1_x:readdata -> mm_interconnect_0:explosion1_x_s1_readdata
	wire   [1:0] mm_interconnect_0_explosion1_x_s1_address;                   // mm_interconnect_0:explosion1_x_s1_address -> explosion1_x:address
	wire         mm_interconnect_0_explosion1_x_s1_write;                     // mm_interconnect_0:explosion1_x_s1_write -> explosion1_x:write_n
	wire  [31:0] mm_interconnect_0_explosion1_x_s1_writedata;                 // mm_interconnect_0:explosion1_x_s1_writedata -> explosion1_x:writedata
	wire         mm_interconnect_0_explosion1_y_s1_chipselect;                // mm_interconnect_0:explosion1_y_s1_chipselect -> explosion1_y:chipselect
	wire  [31:0] mm_interconnect_0_explosion1_y_s1_readdata;                  // explosion1_y:readdata -> mm_interconnect_0:explosion1_y_s1_readdata
	wire   [1:0] mm_interconnect_0_explosion1_y_s1_address;                   // mm_interconnect_0:explosion1_y_s1_address -> explosion1_y:address
	wire         mm_interconnect_0_explosion1_y_s1_write;                     // mm_interconnect_0:explosion1_y_s1_write -> explosion1_y:write_n
	wire  [31:0] mm_interconnect_0_explosion1_y_s1_writedata;                 // mm_interconnect_0:explosion1_y_s1_writedata -> explosion1_y:writedata
	wire         mm_interconnect_0_explosion2_en_s1_chipselect;               // mm_interconnect_0:explosion2_en_s1_chipselect -> explosion2_en:chipselect
	wire  [31:0] mm_interconnect_0_explosion2_en_s1_readdata;                 // explosion2_en:readdata -> mm_interconnect_0:explosion2_en_s1_readdata
	wire   [1:0] mm_interconnect_0_explosion2_en_s1_address;                  // mm_interconnect_0:explosion2_en_s1_address -> explosion2_en:address
	wire         mm_interconnect_0_explosion2_en_s1_write;                    // mm_interconnect_0:explosion2_en_s1_write -> explosion2_en:write_n
	wire  [31:0] mm_interconnect_0_explosion2_en_s1_writedata;                // mm_interconnect_0:explosion2_en_s1_writedata -> explosion2_en:writedata
	wire         mm_interconnect_0_explosion2_x_s1_chipselect;                // mm_interconnect_0:explosion2_x_s1_chipselect -> explosion2_x:chipselect
	wire  [31:0] mm_interconnect_0_explosion2_x_s1_readdata;                  // explosion2_x:readdata -> mm_interconnect_0:explosion2_x_s1_readdata
	wire   [1:0] mm_interconnect_0_explosion2_x_s1_address;                   // mm_interconnect_0:explosion2_x_s1_address -> explosion2_x:address
	wire         mm_interconnect_0_explosion2_x_s1_write;                     // mm_interconnect_0:explosion2_x_s1_write -> explosion2_x:write_n
	wire  [31:0] mm_interconnect_0_explosion2_x_s1_writedata;                 // mm_interconnect_0:explosion2_x_s1_writedata -> explosion2_x:writedata
	wire         mm_interconnect_0_explosion2_y_s1_chipselect;                // mm_interconnect_0:explosion2_y_s1_chipselect -> explosion2_y:chipselect
	wire  [31:0] mm_interconnect_0_explosion2_y_s1_readdata;                  // explosion2_y:readdata -> mm_interconnect_0:explosion2_y_s1_readdata
	wire   [1:0] mm_interconnect_0_explosion2_y_s1_address;                   // mm_interconnect_0:explosion2_y_s1_address -> explosion2_y:address
	wire         mm_interconnect_0_explosion2_y_s1_write;                     // mm_interconnect_0:explosion2_y_s1_write -> explosion2_y:write_n
	wire  [31:0] mm_interconnect_0_explosion2_y_s1_writedata;                 // mm_interconnect_0:explosion2_y_s1_writedata -> explosion2_y:writedata
	wire         mm_interconnect_0_explosion3_en_s1_chipselect;               // mm_interconnect_0:explosion3_en_s1_chipselect -> explosion3_en:chipselect
	wire  [31:0] mm_interconnect_0_explosion3_en_s1_readdata;                 // explosion3_en:readdata -> mm_interconnect_0:explosion3_en_s1_readdata
	wire   [1:0] mm_interconnect_0_explosion3_en_s1_address;                  // mm_interconnect_0:explosion3_en_s1_address -> explosion3_en:address
	wire         mm_interconnect_0_explosion3_en_s1_write;                    // mm_interconnect_0:explosion3_en_s1_write -> explosion3_en:write_n
	wire  [31:0] mm_interconnect_0_explosion3_en_s1_writedata;                // mm_interconnect_0:explosion3_en_s1_writedata -> explosion3_en:writedata
	wire         mm_interconnect_0_explosion3_x_s1_chipselect;                // mm_interconnect_0:explosion3_x_s1_chipselect -> explosion3_x:chipselect
	wire  [31:0] mm_interconnect_0_explosion3_x_s1_readdata;                  // explosion3_x:readdata -> mm_interconnect_0:explosion3_x_s1_readdata
	wire   [1:0] mm_interconnect_0_explosion3_x_s1_address;                   // mm_interconnect_0:explosion3_x_s1_address -> explosion3_x:address
	wire         mm_interconnect_0_explosion3_x_s1_write;                     // mm_interconnect_0:explosion3_x_s1_write -> explosion3_x:write_n
	wire  [31:0] mm_interconnect_0_explosion3_x_s1_writedata;                 // mm_interconnect_0:explosion3_x_s1_writedata -> explosion3_x:writedata
	wire         mm_interconnect_0_explosion3_y_s1_chipselect;                // mm_interconnect_0:explosion3_y_s1_chipselect -> explosion3_y:chipselect
	wire  [31:0] mm_interconnect_0_explosion3_y_s1_readdata;                  // explosion3_y:readdata -> mm_interconnect_0:explosion3_y_s1_readdata
	wire   [1:0] mm_interconnect_0_explosion3_y_s1_address;                   // mm_interconnect_0:explosion3_y_s1_address -> explosion3_y:address
	wire         mm_interconnect_0_explosion3_y_s1_write;                     // mm_interconnect_0:explosion3_y_s1_write -> explosion3_y:write_n
	wire  [31:0] mm_interconnect_0_explosion3_y_s1_writedata;                 // mm_interconnect_0:explosion3_y_s1_writedata -> explosion3_y:writedata
	wire         mm_interconnect_0_bullet1_en_s1_chipselect;                  // mm_interconnect_0:bullet1_en_s1_chipselect -> bullet1_en:chipselect
	wire  [31:0] mm_interconnect_0_bullet1_en_s1_readdata;                    // bullet1_en:readdata -> mm_interconnect_0:bullet1_en_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet1_en_s1_address;                     // mm_interconnect_0:bullet1_en_s1_address -> bullet1_en:address
	wire         mm_interconnect_0_bullet1_en_s1_write;                       // mm_interconnect_0:bullet1_en_s1_write -> bullet1_en:write_n
	wire  [31:0] mm_interconnect_0_bullet1_en_s1_writedata;                   // mm_interconnect_0:bullet1_en_s1_writedata -> bullet1_en:writedata
	wire         mm_interconnect_0_bullet1_x_s1_chipselect;                   // mm_interconnect_0:bullet1_x_s1_chipselect -> bullet1_x:chipselect
	wire  [31:0] mm_interconnect_0_bullet1_x_s1_readdata;                     // bullet1_x:readdata -> mm_interconnect_0:bullet1_x_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet1_x_s1_address;                      // mm_interconnect_0:bullet1_x_s1_address -> bullet1_x:address
	wire         mm_interconnect_0_bullet1_x_s1_write;                        // mm_interconnect_0:bullet1_x_s1_write -> bullet1_x:write_n
	wire  [31:0] mm_interconnect_0_bullet1_x_s1_writedata;                    // mm_interconnect_0:bullet1_x_s1_writedata -> bullet1_x:writedata
	wire         mm_interconnect_0_bullet1_y_s1_chipselect;                   // mm_interconnect_0:bullet1_y_s1_chipselect -> bullet1_y:chipselect
	wire  [31:0] mm_interconnect_0_bullet1_y_s1_readdata;                     // bullet1_y:readdata -> mm_interconnect_0:bullet1_y_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet1_y_s1_address;                      // mm_interconnect_0:bullet1_y_s1_address -> bullet1_y:address
	wire         mm_interconnect_0_bullet1_y_s1_write;                        // mm_interconnect_0:bullet1_y_s1_write -> bullet1_y:write_n
	wire  [31:0] mm_interconnect_0_bullet1_y_s1_writedata;                    // mm_interconnect_0:bullet1_y_s1_writedata -> bullet1_y:writedata
	wire         mm_interconnect_0_bullet2_en_s1_chipselect;                  // mm_interconnect_0:bullet2_en_s1_chipselect -> bullet2_en:chipselect
	wire  [31:0] mm_interconnect_0_bullet2_en_s1_readdata;                    // bullet2_en:readdata -> mm_interconnect_0:bullet2_en_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet2_en_s1_address;                     // mm_interconnect_0:bullet2_en_s1_address -> bullet2_en:address
	wire         mm_interconnect_0_bullet2_en_s1_write;                       // mm_interconnect_0:bullet2_en_s1_write -> bullet2_en:write_n
	wire  [31:0] mm_interconnect_0_bullet2_en_s1_writedata;                   // mm_interconnect_0:bullet2_en_s1_writedata -> bullet2_en:writedata
	wire         mm_interconnect_0_bullet2_x_s1_chipselect;                   // mm_interconnect_0:bullet2_x_s1_chipselect -> bullet2_x:chipselect
	wire  [31:0] mm_interconnect_0_bullet2_x_s1_readdata;                     // bullet2_x:readdata -> mm_interconnect_0:bullet2_x_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet2_x_s1_address;                      // mm_interconnect_0:bullet2_x_s1_address -> bullet2_x:address
	wire         mm_interconnect_0_bullet2_x_s1_write;                        // mm_interconnect_0:bullet2_x_s1_write -> bullet2_x:write_n
	wire  [31:0] mm_interconnect_0_bullet2_x_s1_writedata;                    // mm_interconnect_0:bullet2_x_s1_writedata -> bullet2_x:writedata
	wire         mm_interconnect_0_bullet2_y_s1_chipselect;                   // mm_interconnect_0:bullet2_y_s1_chipselect -> bullet2_y:chipselect
	wire  [31:0] mm_interconnect_0_bullet2_y_s1_readdata;                     // bullet2_y:readdata -> mm_interconnect_0:bullet2_y_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet2_y_s1_address;                      // mm_interconnect_0:bullet2_y_s1_address -> bullet2_y:address
	wire         mm_interconnect_0_bullet2_y_s1_write;                        // mm_interconnect_0:bullet2_y_s1_write -> bullet2_y:write_n
	wire  [31:0] mm_interconnect_0_bullet2_y_s1_writedata;                    // mm_interconnect_0:bullet2_y_s1_writedata -> bullet2_y:writedata
	wire         mm_interconnect_0_bullet3_en_s1_chipselect;                  // mm_interconnect_0:bullet3_en_s1_chipselect -> bullet3_en:chipselect
	wire  [31:0] mm_interconnect_0_bullet3_en_s1_readdata;                    // bullet3_en:readdata -> mm_interconnect_0:bullet3_en_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet3_en_s1_address;                     // mm_interconnect_0:bullet3_en_s1_address -> bullet3_en:address
	wire         mm_interconnect_0_bullet3_en_s1_write;                       // mm_interconnect_0:bullet3_en_s1_write -> bullet3_en:write_n
	wire  [31:0] mm_interconnect_0_bullet3_en_s1_writedata;                   // mm_interconnect_0:bullet3_en_s1_writedata -> bullet3_en:writedata
	wire         mm_interconnect_0_bullet3_x_s1_chipselect;                   // mm_interconnect_0:bullet3_x_s1_chipselect -> bullet3_x:chipselect
	wire  [31:0] mm_interconnect_0_bullet3_x_s1_readdata;                     // bullet3_x:readdata -> mm_interconnect_0:bullet3_x_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet3_x_s1_address;                      // mm_interconnect_0:bullet3_x_s1_address -> bullet3_x:address
	wire         mm_interconnect_0_bullet3_x_s1_write;                        // mm_interconnect_0:bullet3_x_s1_write -> bullet3_x:write_n
	wire  [31:0] mm_interconnect_0_bullet3_x_s1_writedata;                    // mm_interconnect_0:bullet3_x_s1_writedata -> bullet3_x:writedata
	wire         mm_interconnect_0_bullet3_y_s1_chipselect;                   // mm_interconnect_0:bullet3_y_s1_chipselect -> bullet3_y:chipselect
	wire  [31:0] mm_interconnect_0_bullet3_y_s1_readdata;                     // bullet3_y:readdata -> mm_interconnect_0:bullet3_y_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet3_y_s1_address;                      // mm_interconnect_0:bullet3_y_s1_address -> bullet3_y:address
	wire         mm_interconnect_0_bullet3_y_s1_write;                        // mm_interconnect_0:bullet3_y_s1_write -> bullet3_y:write_n
	wire  [31:0] mm_interconnect_0_bullet3_y_s1_writedata;                    // mm_interconnect_0:bullet3_y_s1_writedata -> bullet3_y:writedata
	wire         mm_interconnect_0_health_s1_chipselect;                      // mm_interconnect_0:health_s1_chipselect -> health:chipselect
	wire  [31:0] mm_interconnect_0_health_s1_readdata;                        // health:readdata -> mm_interconnect_0:health_s1_readdata
	wire   [1:0] mm_interconnect_0_health_s1_address;                         // mm_interconnect_0:health_s1_address -> health:address
	wire         mm_interconnect_0_health_s1_write;                           // mm_interconnect_0:health_s1_write -> health:write_n
	wire  [31:0] mm_interconnect_0_health_s1_writedata;                       // mm_interconnect_0:health_s1_writedata -> health:writedata
	wire         mm_interconnect_0_title_en_s1_chipselect;                    // mm_interconnect_0:title_en_s1_chipselect -> title_en:chipselect
	wire  [31:0] mm_interconnect_0_title_en_s1_readdata;                      // title_en:readdata -> mm_interconnect_0:title_en_s1_readdata
	wire   [1:0] mm_interconnect_0_title_en_s1_address;                       // mm_interconnect_0:title_en_s1_address -> title_en:address
	wire         mm_interconnect_0_title_en_s1_write;                         // mm_interconnect_0:title_en_s1_write -> title_en:write_n
	wire  [31:0] mm_interconnect_0_title_en_s1_writedata;                     // mm_interconnect_0:title_en_s1_writedata -> title_en:writedata
	wire         mm_interconnect_0_loss_en_s1_chipselect;                     // mm_interconnect_0:loss_en_s1_chipselect -> loss_en:chipselect
	wire  [31:0] mm_interconnect_0_loss_en_s1_readdata;                       // loss_en:readdata -> mm_interconnect_0:loss_en_s1_readdata
	wire   [1:0] mm_interconnect_0_loss_en_s1_address;                        // mm_interconnect_0:loss_en_s1_address -> loss_en:address
	wire         mm_interconnect_0_loss_en_s1_write;                          // mm_interconnect_0:loss_en_s1_write -> loss_en:write_n
	wire  [31:0] mm_interconnect_0_loss_en_s1_writedata;                      // mm_interconnect_0:loss_en_s1_writedata -> loss_en:writedata
	wire         mm_interconnect_0_win_en_s1_chipselect;                      // mm_interconnect_0:win_en_s1_chipselect -> win_en:chipselect
	wire  [31:0] mm_interconnect_0_win_en_s1_readdata;                        // win_en:readdata -> mm_interconnect_0:win_en_s1_readdata
	wire   [1:0] mm_interconnect_0_win_en_s1_address;                         // mm_interconnect_0:win_en_s1_address -> win_en:address
	wire         mm_interconnect_0_win_en_s1_write;                           // mm_interconnect_0:win_en_s1_write -> win_en:write_n
	wire  [31:0] mm_interconnect_0_win_en_s1_writedata;                       // mm_interconnect_0:win_en_s1_writedata -> win_en:writedata
	wire         mm_interconnect_0_samus_dir_s1_chipselect;                   // mm_interconnect_0:samus_dir_s1_chipselect -> samus_dir:chipselect
	wire  [31:0] mm_interconnect_0_samus_dir_s1_readdata;                     // samus_dir:readdata -> mm_interconnect_0:samus_dir_s1_readdata
	wire   [1:0] mm_interconnect_0_samus_dir_s1_address;                      // mm_interconnect_0:samus_dir_s1_address -> samus_dir:address
	wire         mm_interconnect_0_samus_dir_s1_write;                        // mm_interconnect_0:samus_dir_s1_write -> samus_dir:write_n
	wire  [31:0] mm_interconnect_0_samus_dir_s1_writedata;                    // mm_interconnect_0:samus_dir_s1_writedata -> samus_dir:writedata
	wire         mm_interconnect_0_scene_sel_s1_chipselect;                   // mm_interconnect_0:scene_sel_s1_chipselect -> scene_sel:chipselect
	wire  [31:0] mm_interconnect_0_scene_sel_s1_readdata;                     // scene_sel:readdata -> mm_interconnect_0:scene_sel_s1_readdata
	wire   [1:0] mm_interconnect_0_scene_sel_s1_address;                      // mm_interconnect_0:scene_sel_s1_address -> scene_sel:address
	wire         mm_interconnect_0_scene_sel_s1_write;                        // mm_interconnect_0:scene_sel_s1_write -> scene_sel:write_n
	wire  [31:0] mm_interconnect_0_scene_sel_s1_writedata;                    // mm_interconnect_0:scene_sel_s1_writedata -> scene_sel:writedata
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_qsys_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_qsys_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [bullet1_en:reset_n, bullet1_x:reset_n, bullet1_y:reset_n, bullet2_en:reset_n, bullet2_x:reset_n, bullet2_y:reset_n, bullet3_en:reset_n, bullet3_x:reset_n, bullet3_y:reset_n, explosion1_en:reset_n, explosion1_x:reset_n, explosion1_y:reset_n, explosion2_en:reset_n, explosion2_x:reset_n, explosion2_y:reset_n, explosion3_en:reset_n, explosion3_x:reset_n, explosion3_y:reset_n, health:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, key:reset_n, keycode:reset_n, loss_en:reset_n, mm_interconnect_0:nios2_qsys_0_reset_reset_bridge_in_reset_reset, monster1_en:reset_n, monster1_x:reset_n, monster1_y:reset_n, monster2_en:reset_n, monster2_x:reset_n, monster2_y:reset_n, monster3_en:reset_n, monster3_x:reset_n, monster3_y:reset_n, nios2_qsys_0:reset_n, onchip_memory2_0:reset, otg_hpi_address:reset_n, otg_hpi_cs:reset_n, otg_hpi_data:reset_n, otg_hpi_r:reset_n, otg_hpi_w:reset_n, rst_translator:in_reset, samus_dir:reset_n, samus_en:reset_n, samus_jump:reset_n, samus_walk:reset_n, samus_x:reset_n, samus_y:reset_n, scene_sel:reset_n, sdram_pll:reset, sysid_qsys_0:reset_n, title_en:reset_n, win_en:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [nios2_qsys_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_qsys_0_debug_reset_request_reset;                      // nios2_qsys_0:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [mm_interconnect_0:sdram_reset_reset_bridge_in_reset_reset, sdram:reset_n]

	nios_system_bullet1_en bullet1_en (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_bullet1_en_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet1_en_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet1_en_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet1_en_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet1_en_s1_readdata),   //                    .readdata
		.out_port   (bullet1_en_export)                           // external_connection.export
	);

	nios_system_bullet1_x bullet1_x (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_bullet1_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet1_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet1_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet1_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet1_x_s1_readdata),   //                    .readdata
		.out_port   (bullet1_x_export)                           // external_connection.export
	);

	nios_system_bullet1_x bullet1_y (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_bullet1_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet1_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet1_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet1_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet1_y_s1_readdata),   //                    .readdata
		.out_port   (bullet1_y_export)                           // external_connection.export
	);

	nios_system_bullet1_en bullet2_en (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_bullet2_en_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet2_en_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet2_en_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet2_en_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet2_en_s1_readdata),   //                    .readdata
		.out_port   (bullet2_en_export)                           // external_connection.export
	);

	nios_system_bullet1_x bullet2_x (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_bullet2_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet2_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet2_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet2_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet2_x_s1_readdata),   //                    .readdata
		.out_port   (bullet2_x_export)                           // external_connection.export
	);

	nios_system_bullet1_x bullet2_y (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_bullet2_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet2_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet2_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet2_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet2_y_s1_readdata),   //                    .readdata
		.out_port   (bullet2_y_export)                           // external_connection.export
	);

	nios_system_bullet1_en bullet3_en (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_bullet3_en_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet3_en_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet3_en_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet3_en_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet3_en_s1_readdata),   //                    .readdata
		.out_port   (bullet3_en_export)                           // external_connection.export
	);

	nios_system_bullet1_x bullet3_x (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_bullet3_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet3_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet3_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet3_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet3_x_s1_readdata),   //                    .readdata
		.out_port   (bullet3_x_export)                           // external_connection.export
	);

	nios_system_bullet1_x bullet3_y (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_bullet3_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet3_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet3_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet3_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet3_y_s1_readdata),   //                    .readdata
		.out_port   (bullet3_y_export)                           // external_connection.export
	);

	nios_system_bullet1_en explosion1_en (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_explosion1_en_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_explosion1_en_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_explosion1_en_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_explosion1_en_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_explosion1_en_s1_readdata),   //                    .readdata
		.out_port   (explosion1_en_export)                           // external_connection.export
	);

	nios_system_bullet1_x explosion1_x (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_explosion1_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_explosion1_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_explosion1_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_explosion1_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_explosion1_x_s1_readdata),   //                    .readdata
		.out_port   (explosion1_x_export)                           // external_connection.export
	);

	nios_system_bullet1_x explosion1_y (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_explosion1_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_explosion1_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_explosion1_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_explosion1_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_explosion1_y_s1_readdata),   //                    .readdata
		.out_port   (explosion1_y_export)                           // external_connection.export
	);

	nios_system_bullet1_en explosion2_en (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_explosion2_en_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_explosion2_en_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_explosion2_en_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_explosion2_en_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_explosion2_en_s1_readdata),   //                    .readdata
		.out_port   (explosion2_en_export)                           // external_connection.export
	);

	nios_system_bullet1_x explosion2_x (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_explosion2_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_explosion2_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_explosion2_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_explosion2_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_explosion2_x_s1_readdata),   //                    .readdata
		.out_port   (explosion2_x_export)                           // external_connection.export
	);

	nios_system_bullet1_x explosion2_y (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_explosion2_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_explosion2_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_explosion2_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_explosion2_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_explosion2_y_s1_readdata),   //                    .readdata
		.out_port   (explosion2_y_export)                           // external_connection.export
	);

	nios_system_bullet1_en explosion3_en (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_explosion3_en_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_explosion3_en_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_explosion3_en_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_explosion3_en_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_explosion3_en_s1_readdata),   //                    .readdata
		.out_port   (explosion3_en_export)                           // external_connection.export
	);

	nios_system_bullet1_x explosion3_x (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_explosion3_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_explosion3_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_explosion3_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_explosion3_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_explosion3_x_s1_readdata),   //                    .readdata
		.out_port   (explosion3_x_export)                           // external_connection.export
	);

	nios_system_bullet1_x explosion3_y (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_explosion3_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_explosion3_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_explosion3_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_explosion3_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_explosion3_y_s1_readdata),   //                    .readdata
		.out_port   (explosion3_y_export)                           // external_connection.export
	);

	nios_system_health health (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_health_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_health_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_health_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_health_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_health_s1_readdata),   //                    .readdata
		.out_port   (health_export)                           // external_connection.export
	);

	nios_system_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	nios_system_key key (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_key_s1_readdata),   //                    .readdata
		.in_port    (key_export)                           // external_connection.export
	);

	nios_system_keycode keycode (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_keycode_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_keycode_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_keycode_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_keycode_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_keycode_s1_readdata),   //                    .readdata
		.out_port   (keycode_export)                           // external_connection.export
	);

	nios_system_bullet1_en loss_en (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_loss_en_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_loss_en_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_loss_en_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_loss_en_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_loss_en_s1_readdata),   //                    .readdata
		.out_port   (loss_en_export)                           // external_connection.export
	);

	nios_system_bullet1_en monster1_en (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_monster1_en_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_monster1_en_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_monster1_en_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_monster1_en_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_monster1_en_s1_readdata),   //                    .readdata
		.out_port   (monster1_en_export)                           // external_connection.export
	);

	nios_system_bullet1_x monster1_x (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_monster1_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_monster1_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_monster1_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_monster1_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_monster1_x_s1_readdata),   //                    .readdata
		.out_port   (monster1_x_export)                           // external_connection.export
	);

	nios_system_bullet1_x monster1_y (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_monster1_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_monster1_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_monster1_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_monster1_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_monster1_y_s1_readdata),   //                    .readdata
		.out_port   (monster1_y_export)                           // external_connection.export
	);

	nios_system_bullet1_en monster2_en (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_monster2_en_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_monster2_en_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_monster2_en_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_monster2_en_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_monster2_en_s1_readdata),   //                    .readdata
		.out_port   (monster2_en_export)                           // external_connection.export
	);

	nios_system_bullet1_x monster2_x (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_monster2_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_monster2_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_monster2_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_monster2_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_monster2_x_s1_readdata),   //                    .readdata
		.out_port   (monster2_x_export)                           // external_connection.export
	);

	nios_system_bullet1_x monster2_y (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_monster2_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_monster2_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_monster2_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_monster2_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_monster2_y_s1_readdata),   //                    .readdata
		.out_port   (monster2_y_export)                           // external_connection.export
	);

	nios_system_bullet1_en monster3_en (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_monster3_en_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_monster3_en_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_monster3_en_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_monster3_en_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_monster3_en_s1_readdata),   //                    .readdata
		.out_port   (monster3_en_export)                           // external_connection.export
	);

	nios_system_bullet1_x monster3_x (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_monster3_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_monster3_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_monster3_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_monster3_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_monster3_x_s1_readdata),   //                    .readdata
		.out_port   (monster3_x_export)                           // external_connection.export
	);

	nios_system_bullet1_x monster3_y (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_monster3_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_monster3_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_monster3_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_monster3_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_monster3_y_s1_readdata),   //                    .readdata
		.out_port   (monster3_y_export)                           // external_connection.export
	);

	nios_system_nios2_qsys_0 nios2_qsys_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_qsys_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_qsys_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_qsys_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_qsys_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_qsys_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_qsys_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_qsys_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_qsys_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_qsys_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_qsys_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_qsys_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_qsys_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_qsys_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	nios_system_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                //       .reset_req
	);

	nios_system_health otg_hpi_address (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_address_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_address_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_address_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_address_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_address_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_address_export)                           // external_connection.export
	);

	nios_system_bullet1_en otg_hpi_cs (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_cs_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_cs_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_cs_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_cs_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_cs_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_cs_export)                           // external_connection.export
	);

	nios_system_otg_hpi_data otg_hpi_data (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_data_s1_readdata),   //                    .readdata
		.in_port    (otg_hpi_data_in_port),                         // external_connection.export
		.out_port   (otg_hpi_data_out_port)                         //                    .export
	);

	nios_system_bullet1_en otg_hpi_r (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_r_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_r_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_r_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_r_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_r_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_r_export)                           // external_connection.export
	);

	nios_system_bullet1_en otg_hpi_w (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_w_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_w_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_w_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_w_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_w_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_w_export)                           // external_connection.export
	);

	nios_system_bullet1_en samus_dir (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_samus_dir_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_samus_dir_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_samus_dir_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_samus_dir_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_samus_dir_s1_readdata),   //                    .readdata
		.out_port   (samus_dir_export)                           // external_connection.export
	);

	nios_system_bullet1_en samus_en (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_samus_en_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_samus_en_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_samus_en_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_samus_en_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_samus_en_s1_readdata),   //                    .readdata
		.out_port   (samus_en_export)                           // external_connection.export
	);

	nios_system_bullet1_en samus_jump (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_samus_jump_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_samus_jump_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_samus_jump_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_samus_jump_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_samus_jump_s1_readdata),   //                    .readdata
		.out_port   (samus_jump_export)                           // external_connection.export
	);

	nios_system_bullet1_en samus_walk (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_samus_walk_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_samus_walk_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_samus_walk_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_samus_walk_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_samus_walk_s1_readdata),   //                    .readdata
		.out_port   (samus_walk_export)                           // external_connection.export
	);

	nios_system_bullet1_x samus_x (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_samus_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_samus_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_samus_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_samus_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_samus_x_s1_readdata),   //                    .readdata
		.out_port   (samus_x_export)                           // external_connection.export
	);

	nios_system_bullet1_x samus_y (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_samus_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_samus_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_samus_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_samus_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_samus_y_s1_readdata),   //                    .readdata
		.out_port   (samus_y_export)                           // external_connection.export
	);

	nios_system_scene_sel scene_sel (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_scene_sel_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_scene_sel_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_scene_sel_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_scene_sel_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_scene_sel_s1_readdata),   //                    .readdata
		.out_port   (scene_sel_export)                           // external_connection.export
	);

	nios_system_sdram sdram (
		.clk            (sdram_pll_c0_clk),                         //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	nios_system_sdram_pll sdram_pll (
		.clk       (clk_clk),                                         //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset),                  // inclk_interface_reset.reset
		.read      (mm_interconnect_0_sdram_pll_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_sdram_pll_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_sdram_pll_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_sdram_pll_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_sdram_pll_pll_slave_writedata), //                      .writedata
		.c0        (sdram_pll_c0_clk),                                //                    c0.clk
		.c1        (sdram_clk_clk),                                   //                    c1.clk
		.areset    (),                                                //        areset_conduit.export
		.locked    (),                                                //        locked_conduit.export
		.phasedone ()                                                 //     phasedone_conduit.export
	);

	nios_system_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	nios_system_bullet1_en title_en (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_title_en_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_title_en_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_title_en_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_title_en_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_title_en_s1_readdata),   //                    .readdata
		.out_port   (title_en_export)                           // external_connection.export
	);

	nios_system_bullet1_en win_en (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_win_en_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_win_en_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_win_en_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_win_en_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_win_en_s1_readdata),   //                    .readdata
		.out_port   (win_en_export)                           // external_connection.export
	);

	nios_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                     //                                clk_0_clk.clk
		.sdram_pll_c0_clk                               (sdram_pll_c0_clk),                                            //                             sdram_pll_c0.clk
		.nios2_qsys_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // nios2_qsys_0_reset_reset_bridge_in_reset.reset
		.sdram_reset_reset_bridge_in_reset_reset        (rst_controller_001_reset_out_reset),                          //        sdram_reset_reset_bridge_in_reset.reset
		.nios2_qsys_0_data_master_address               (nios2_qsys_0_data_master_address),                            //                 nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest           (nios2_qsys_0_data_master_waitrequest),                        //                                         .waitrequest
		.nios2_qsys_0_data_master_byteenable            (nios2_qsys_0_data_master_byteenable),                         //                                         .byteenable
		.nios2_qsys_0_data_master_read                  (nios2_qsys_0_data_master_read),                               //                                         .read
		.nios2_qsys_0_data_master_readdata              (nios2_qsys_0_data_master_readdata),                           //                                         .readdata
		.nios2_qsys_0_data_master_write                 (nios2_qsys_0_data_master_write),                              //                                         .write
		.nios2_qsys_0_data_master_writedata             (nios2_qsys_0_data_master_writedata),                          //                                         .writedata
		.nios2_qsys_0_data_master_debugaccess           (nios2_qsys_0_data_master_debugaccess),                        //                                         .debugaccess
		.nios2_qsys_0_instruction_master_address        (nios2_qsys_0_instruction_master_address),                     //          nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest    (nios2_qsys_0_instruction_master_waitrequest),                 //                                         .waitrequest
		.nios2_qsys_0_instruction_master_read           (nios2_qsys_0_instruction_master_read),                        //                                         .read
		.nios2_qsys_0_instruction_master_readdata       (nios2_qsys_0_instruction_master_readdata),                    //                                         .readdata
		.bullet1_en_s1_address                          (mm_interconnect_0_bullet1_en_s1_address),                     //                            bullet1_en_s1.address
		.bullet1_en_s1_write                            (mm_interconnect_0_bullet1_en_s1_write),                       //                                         .write
		.bullet1_en_s1_readdata                         (mm_interconnect_0_bullet1_en_s1_readdata),                    //                                         .readdata
		.bullet1_en_s1_writedata                        (mm_interconnect_0_bullet1_en_s1_writedata),                   //                                         .writedata
		.bullet1_en_s1_chipselect                       (mm_interconnect_0_bullet1_en_s1_chipselect),                  //                                         .chipselect
		.bullet1_x_s1_address                           (mm_interconnect_0_bullet1_x_s1_address),                      //                             bullet1_x_s1.address
		.bullet1_x_s1_write                             (mm_interconnect_0_bullet1_x_s1_write),                        //                                         .write
		.bullet1_x_s1_readdata                          (mm_interconnect_0_bullet1_x_s1_readdata),                     //                                         .readdata
		.bullet1_x_s1_writedata                         (mm_interconnect_0_bullet1_x_s1_writedata),                    //                                         .writedata
		.bullet1_x_s1_chipselect                        (mm_interconnect_0_bullet1_x_s1_chipselect),                   //                                         .chipselect
		.bullet1_y_s1_address                           (mm_interconnect_0_bullet1_y_s1_address),                      //                             bullet1_y_s1.address
		.bullet1_y_s1_write                             (mm_interconnect_0_bullet1_y_s1_write),                        //                                         .write
		.bullet1_y_s1_readdata                          (mm_interconnect_0_bullet1_y_s1_readdata),                     //                                         .readdata
		.bullet1_y_s1_writedata                         (mm_interconnect_0_bullet1_y_s1_writedata),                    //                                         .writedata
		.bullet1_y_s1_chipselect                        (mm_interconnect_0_bullet1_y_s1_chipselect),                   //                                         .chipselect
		.bullet2_en_s1_address                          (mm_interconnect_0_bullet2_en_s1_address),                     //                            bullet2_en_s1.address
		.bullet2_en_s1_write                            (mm_interconnect_0_bullet2_en_s1_write),                       //                                         .write
		.bullet2_en_s1_readdata                         (mm_interconnect_0_bullet2_en_s1_readdata),                    //                                         .readdata
		.bullet2_en_s1_writedata                        (mm_interconnect_0_bullet2_en_s1_writedata),                   //                                         .writedata
		.bullet2_en_s1_chipselect                       (mm_interconnect_0_bullet2_en_s1_chipselect),                  //                                         .chipselect
		.bullet2_x_s1_address                           (mm_interconnect_0_bullet2_x_s1_address),                      //                             bullet2_x_s1.address
		.bullet2_x_s1_write                             (mm_interconnect_0_bullet2_x_s1_write),                        //                                         .write
		.bullet2_x_s1_readdata                          (mm_interconnect_0_bullet2_x_s1_readdata),                     //                                         .readdata
		.bullet2_x_s1_writedata                         (mm_interconnect_0_bullet2_x_s1_writedata),                    //                                         .writedata
		.bullet2_x_s1_chipselect                        (mm_interconnect_0_bullet2_x_s1_chipselect),                   //                                         .chipselect
		.bullet2_y_s1_address                           (mm_interconnect_0_bullet2_y_s1_address),                      //                             bullet2_y_s1.address
		.bullet2_y_s1_write                             (mm_interconnect_0_bullet2_y_s1_write),                        //                                         .write
		.bullet2_y_s1_readdata                          (mm_interconnect_0_bullet2_y_s1_readdata),                     //                                         .readdata
		.bullet2_y_s1_writedata                         (mm_interconnect_0_bullet2_y_s1_writedata),                    //                                         .writedata
		.bullet2_y_s1_chipselect                        (mm_interconnect_0_bullet2_y_s1_chipselect),                   //                                         .chipselect
		.bullet3_en_s1_address                          (mm_interconnect_0_bullet3_en_s1_address),                     //                            bullet3_en_s1.address
		.bullet3_en_s1_write                            (mm_interconnect_0_bullet3_en_s1_write),                       //                                         .write
		.bullet3_en_s1_readdata                         (mm_interconnect_0_bullet3_en_s1_readdata),                    //                                         .readdata
		.bullet3_en_s1_writedata                        (mm_interconnect_0_bullet3_en_s1_writedata),                   //                                         .writedata
		.bullet3_en_s1_chipselect                       (mm_interconnect_0_bullet3_en_s1_chipselect),                  //                                         .chipselect
		.bullet3_x_s1_address                           (mm_interconnect_0_bullet3_x_s1_address),                      //                             bullet3_x_s1.address
		.bullet3_x_s1_write                             (mm_interconnect_0_bullet3_x_s1_write),                        //                                         .write
		.bullet3_x_s1_readdata                          (mm_interconnect_0_bullet3_x_s1_readdata),                     //                                         .readdata
		.bullet3_x_s1_writedata                         (mm_interconnect_0_bullet3_x_s1_writedata),                    //                                         .writedata
		.bullet3_x_s1_chipselect                        (mm_interconnect_0_bullet3_x_s1_chipselect),                   //                                         .chipselect
		.bullet3_y_s1_address                           (mm_interconnect_0_bullet3_y_s1_address),                      //                             bullet3_y_s1.address
		.bullet3_y_s1_write                             (mm_interconnect_0_bullet3_y_s1_write),                        //                                         .write
		.bullet3_y_s1_readdata                          (mm_interconnect_0_bullet3_y_s1_readdata),                     //                                         .readdata
		.bullet3_y_s1_writedata                         (mm_interconnect_0_bullet3_y_s1_writedata),                    //                                         .writedata
		.bullet3_y_s1_chipselect                        (mm_interconnect_0_bullet3_y_s1_chipselect),                   //                                         .chipselect
		.explosion1_en_s1_address                       (mm_interconnect_0_explosion1_en_s1_address),                  //                         explosion1_en_s1.address
		.explosion1_en_s1_write                         (mm_interconnect_0_explosion1_en_s1_write),                    //                                         .write
		.explosion1_en_s1_readdata                      (mm_interconnect_0_explosion1_en_s1_readdata),                 //                                         .readdata
		.explosion1_en_s1_writedata                     (mm_interconnect_0_explosion1_en_s1_writedata),                //                                         .writedata
		.explosion1_en_s1_chipselect                    (mm_interconnect_0_explosion1_en_s1_chipselect),               //                                         .chipselect
		.explosion1_x_s1_address                        (mm_interconnect_0_explosion1_x_s1_address),                   //                          explosion1_x_s1.address
		.explosion1_x_s1_write                          (mm_interconnect_0_explosion1_x_s1_write),                     //                                         .write
		.explosion1_x_s1_readdata                       (mm_interconnect_0_explosion1_x_s1_readdata),                  //                                         .readdata
		.explosion1_x_s1_writedata                      (mm_interconnect_0_explosion1_x_s1_writedata),                 //                                         .writedata
		.explosion1_x_s1_chipselect                     (mm_interconnect_0_explosion1_x_s1_chipselect),                //                                         .chipselect
		.explosion1_y_s1_address                        (mm_interconnect_0_explosion1_y_s1_address),                   //                          explosion1_y_s1.address
		.explosion1_y_s1_write                          (mm_interconnect_0_explosion1_y_s1_write),                     //                                         .write
		.explosion1_y_s1_readdata                       (mm_interconnect_0_explosion1_y_s1_readdata),                  //                                         .readdata
		.explosion1_y_s1_writedata                      (mm_interconnect_0_explosion1_y_s1_writedata),                 //                                         .writedata
		.explosion1_y_s1_chipselect                     (mm_interconnect_0_explosion1_y_s1_chipselect),                //                                         .chipselect
		.explosion2_en_s1_address                       (mm_interconnect_0_explosion2_en_s1_address),                  //                         explosion2_en_s1.address
		.explosion2_en_s1_write                         (mm_interconnect_0_explosion2_en_s1_write),                    //                                         .write
		.explosion2_en_s1_readdata                      (mm_interconnect_0_explosion2_en_s1_readdata),                 //                                         .readdata
		.explosion2_en_s1_writedata                     (mm_interconnect_0_explosion2_en_s1_writedata),                //                                         .writedata
		.explosion2_en_s1_chipselect                    (mm_interconnect_0_explosion2_en_s1_chipselect),               //                                         .chipselect
		.explosion2_x_s1_address                        (mm_interconnect_0_explosion2_x_s1_address),                   //                          explosion2_x_s1.address
		.explosion2_x_s1_write                          (mm_interconnect_0_explosion2_x_s1_write),                     //                                         .write
		.explosion2_x_s1_readdata                       (mm_interconnect_0_explosion2_x_s1_readdata),                  //                                         .readdata
		.explosion2_x_s1_writedata                      (mm_interconnect_0_explosion2_x_s1_writedata),                 //                                         .writedata
		.explosion2_x_s1_chipselect                     (mm_interconnect_0_explosion2_x_s1_chipselect),                //                                         .chipselect
		.explosion2_y_s1_address                        (mm_interconnect_0_explosion2_y_s1_address),                   //                          explosion2_y_s1.address
		.explosion2_y_s1_write                          (mm_interconnect_0_explosion2_y_s1_write),                     //                                         .write
		.explosion2_y_s1_readdata                       (mm_interconnect_0_explosion2_y_s1_readdata),                  //                                         .readdata
		.explosion2_y_s1_writedata                      (mm_interconnect_0_explosion2_y_s1_writedata),                 //                                         .writedata
		.explosion2_y_s1_chipselect                     (mm_interconnect_0_explosion2_y_s1_chipselect),                //                                         .chipselect
		.explosion3_en_s1_address                       (mm_interconnect_0_explosion3_en_s1_address),                  //                         explosion3_en_s1.address
		.explosion3_en_s1_write                         (mm_interconnect_0_explosion3_en_s1_write),                    //                                         .write
		.explosion3_en_s1_readdata                      (mm_interconnect_0_explosion3_en_s1_readdata),                 //                                         .readdata
		.explosion3_en_s1_writedata                     (mm_interconnect_0_explosion3_en_s1_writedata),                //                                         .writedata
		.explosion3_en_s1_chipselect                    (mm_interconnect_0_explosion3_en_s1_chipselect),               //                                         .chipselect
		.explosion3_x_s1_address                        (mm_interconnect_0_explosion3_x_s1_address),                   //                          explosion3_x_s1.address
		.explosion3_x_s1_write                          (mm_interconnect_0_explosion3_x_s1_write),                     //                                         .write
		.explosion3_x_s1_readdata                       (mm_interconnect_0_explosion3_x_s1_readdata),                  //                                         .readdata
		.explosion3_x_s1_writedata                      (mm_interconnect_0_explosion3_x_s1_writedata),                 //                                         .writedata
		.explosion3_x_s1_chipselect                     (mm_interconnect_0_explosion3_x_s1_chipselect),                //                                         .chipselect
		.explosion3_y_s1_address                        (mm_interconnect_0_explosion3_y_s1_address),                   //                          explosion3_y_s1.address
		.explosion3_y_s1_write                          (mm_interconnect_0_explosion3_y_s1_write),                     //                                         .write
		.explosion3_y_s1_readdata                       (mm_interconnect_0_explosion3_y_s1_readdata),                  //                                         .readdata
		.explosion3_y_s1_writedata                      (mm_interconnect_0_explosion3_y_s1_writedata),                 //                                         .writedata
		.explosion3_y_s1_chipselect                     (mm_interconnect_0_explosion3_y_s1_chipselect),                //                                         .chipselect
		.health_s1_address                              (mm_interconnect_0_health_s1_address),                         //                                health_s1.address
		.health_s1_write                                (mm_interconnect_0_health_s1_write),                           //                                         .write
		.health_s1_readdata                             (mm_interconnect_0_health_s1_readdata),                        //                                         .readdata
		.health_s1_writedata                            (mm_interconnect_0_health_s1_writedata),                       //                                         .writedata
		.health_s1_chipselect                           (mm_interconnect_0_health_s1_chipselect),                      //                                         .chipselect
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.key_s1_address                                 (mm_interconnect_0_key_s1_address),                            //                                   key_s1.address
		.key_s1_write                                   (mm_interconnect_0_key_s1_write),                              //                                         .write
		.key_s1_readdata                                (mm_interconnect_0_key_s1_readdata),                           //                                         .readdata
		.key_s1_writedata                               (mm_interconnect_0_key_s1_writedata),                          //                                         .writedata
		.key_s1_chipselect                              (mm_interconnect_0_key_s1_chipselect),                         //                                         .chipselect
		.keycode_s1_address                             (mm_interconnect_0_keycode_s1_address),                        //                               keycode_s1.address
		.keycode_s1_write                               (mm_interconnect_0_keycode_s1_write),                          //                                         .write
		.keycode_s1_readdata                            (mm_interconnect_0_keycode_s1_readdata),                       //                                         .readdata
		.keycode_s1_writedata                           (mm_interconnect_0_keycode_s1_writedata),                      //                                         .writedata
		.keycode_s1_chipselect                          (mm_interconnect_0_keycode_s1_chipselect),                     //                                         .chipselect
		.loss_en_s1_address                             (mm_interconnect_0_loss_en_s1_address),                        //                               loss_en_s1.address
		.loss_en_s1_write                               (mm_interconnect_0_loss_en_s1_write),                          //                                         .write
		.loss_en_s1_readdata                            (mm_interconnect_0_loss_en_s1_readdata),                       //                                         .readdata
		.loss_en_s1_writedata                           (mm_interconnect_0_loss_en_s1_writedata),                      //                                         .writedata
		.loss_en_s1_chipselect                          (mm_interconnect_0_loss_en_s1_chipselect),                     //                                         .chipselect
		.monster1_en_s1_address                         (mm_interconnect_0_monster1_en_s1_address),                    //                           monster1_en_s1.address
		.monster1_en_s1_write                           (mm_interconnect_0_monster1_en_s1_write),                      //                                         .write
		.monster1_en_s1_readdata                        (mm_interconnect_0_monster1_en_s1_readdata),                   //                                         .readdata
		.monster1_en_s1_writedata                       (mm_interconnect_0_monster1_en_s1_writedata),                  //                                         .writedata
		.monster1_en_s1_chipselect                      (mm_interconnect_0_monster1_en_s1_chipselect),                 //                                         .chipselect
		.monster1_x_s1_address                          (mm_interconnect_0_monster1_x_s1_address),                     //                            monster1_x_s1.address
		.monster1_x_s1_write                            (mm_interconnect_0_monster1_x_s1_write),                       //                                         .write
		.monster1_x_s1_readdata                         (mm_interconnect_0_monster1_x_s1_readdata),                    //                                         .readdata
		.monster1_x_s1_writedata                        (mm_interconnect_0_monster1_x_s1_writedata),                   //                                         .writedata
		.monster1_x_s1_chipselect                       (mm_interconnect_0_monster1_x_s1_chipselect),                  //                                         .chipselect
		.monster1_y_s1_address                          (mm_interconnect_0_monster1_y_s1_address),                     //                            monster1_y_s1.address
		.monster1_y_s1_write                            (mm_interconnect_0_monster1_y_s1_write),                       //                                         .write
		.monster1_y_s1_readdata                         (mm_interconnect_0_monster1_y_s1_readdata),                    //                                         .readdata
		.monster1_y_s1_writedata                        (mm_interconnect_0_monster1_y_s1_writedata),                   //                                         .writedata
		.monster1_y_s1_chipselect                       (mm_interconnect_0_monster1_y_s1_chipselect),                  //                                         .chipselect
		.monster2_en_s1_address                         (mm_interconnect_0_monster2_en_s1_address),                    //                           monster2_en_s1.address
		.monster2_en_s1_write                           (mm_interconnect_0_monster2_en_s1_write),                      //                                         .write
		.monster2_en_s1_readdata                        (mm_interconnect_0_monster2_en_s1_readdata),                   //                                         .readdata
		.monster2_en_s1_writedata                       (mm_interconnect_0_monster2_en_s1_writedata),                  //                                         .writedata
		.monster2_en_s1_chipselect                      (mm_interconnect_0_monster2_en_s1_chipselect),                 //                                         .chipselect
		.monster2_x_s1_address                          (mm_interconnect_0_monster2_x_s1_address),                     //                            monster2_x_s1.address
		.monster2_x_s1_write                            (mm_interconnect_0_monster2_x_s1_write),                       //                                         .write
		.monster2_x_s1_readdata                         (mm_interconnect_0_monster2_x_s1_readdata),                    //                                         .readdata
		.monster2_x_s1_writedata                        (mm_interconnect_0_monster2_x_s1_writedata),                   //                                         .writedata
		.monster2_x_s1_chipselect                       (mm_interconnect_0_monster2_x_s1_chipselect),                  //                                         .chipselect
		.monster2_y_s1_address                          (mm_interconnect_0_monster2_y_s1_address),                     //                            monster2_y_s1.address
		.monster2_y_s1_write                            (mm_interconnect_0_monster2_y_s1_write),                       //                                         .write
		.monster2_y_s1_readdata                         (mm_interconnect_0_monster2_y_s1_readdata),                    //                                         .readdata
		.monster2_y_s1_writedata                        (mm_interconnect_0_monster2_y_s1_writedata),                   //                                         .writedata
		.monster2_y_s1_chipselect                       (mm_interconnect_0_monster2_y_s1_chipselect),                  //                                         .chipselect
		.monster3_en_s1_address                         (mm_interconnect_0_monster3_en_s1_address),                    //                           monster3_en_s1.address
		.monster3_en_s1_write                           (mm_interconnect_0_monster3_en_s1_write),                      //                                         .write
		.monster3_en_s1_readdata                        (mm_interconnect_0_monster3_en_s1_readdata),                   //                                         .readdata
		.monster3_en_s1_writedata                       (mm_interconnect_0_monster3_en_s1_writedata),                  //                                         .writedata
		.monster3_en_s1_chipselect                      (mm_interconnect_0_monster3_en_s1_chipselect),                 //                                         .chipselect
		.monster3_x_s1_address                          (mm_interconnect_0_monster3_x_s1_address),                     //                            monster3_x_s1.address
		.monster3_x_s1_write                            (mm_interconnect_0_monster3_x_s1_write),                       //                                         .write
		.monster3_x_s1_readdata                         (mm_interconnect_0_monster3_x_s1_readdata),                    //                                         .readdata
		.monster3_x_s1_writedata                        (mm_interconnect_0_monster3_x_s1_writedata),                   //                                         .writedata
		.monster3_x_s1_chipselect                       (mm_interconnect_0_monster3_x_s1_chipselect),                  //                                         .chipselect
		.monster3_y_s1_address                          (mm_interconnect_0_monster3_y_s1_address),                     //                            monster3_y_s1.address
		.monster3_y_s1_write                            (mm_interconnect_0_monster3_y_s1_write),                       //                                         .write
		.monster3_y_s1_readdata                         (mm_interconnect_0_monster3_y_s1_readdata),                    //                                         .readdata
		.monster3_y_s1_writedata                        (mm_interconnect_0_monster3_y_s1_writedata),                   //                                         .writedata
		.monster3_y_s1_chipselect                       (mm_interconnect_0_monster3_y_s1_chipselect),                  //                                         .chipselect
		.nios2_qsys_0_debug_mem_slave_address           (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_address),      //             nios2_qsys_0_debug_mem_slave.address
		.nios2_qsys_0_debug_mem_slave_write             (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_write),        //                                         .write
		.nios2_qsys_0_debug_mem_slave_read              (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_read),         //                                         .read
		.nios2_qsys_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_readdata),     //                                         .readdata
		.nios2_qsys_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_writedata),    //                                         .writedata
		.nios2_qsys_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_byteenable),   //                                         .byteenable
		.nios2_qsys_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_waitrequest),  //                                         .waitrequest
		.nios2_qsys_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_debugaccess),  //                                         .debugaccess
		.onchip_memory2_0_s1_address                    (mm_interconnect_0_onchip_memory2_0_s1_address),               //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                         .clken
		.otg_hpi_address_s1_address                     (mm_interconnect_0_otg_hpi_address_s1_address),                //                       otg_hpi_address_s1.address
		.otg_hpi_address_s1_write                       (mm_interconnect_0_otg_hpi_address_s1_write),                  //                                         .write
		.otg_hpi_address_s1_readdata                    (mm_interconnect_0_otg_hpi_address_s1_readdata),               //                                         .readdata
		.otg_hpi_address_s1_writedata                   (mm_interconnect_0_otg_hpi_address_s1_writedata),              //                                         .writedata
		.otg_hpi_address_s1_chipselect                  (mm_interconnect_0_otg_hpi_address_s1_chipselect),             //                                         .chipselect
		.otg_hpi_cs_s1_address                          (mm_interconnect_0_otg_hpi_cs_s1_address),                     //                            otg_hpi_cs_s1.address
		.otg_hpi_cs_s1_write                            (mm_interconnect_0_otg_hpi_cs_s1_write),                       //                                         .write
		.otg_hpi_cs_s1_readdata                         (mm_interconnect_0_otg_hpi_cs_s1_readdata),                    //                                         .readdata
		.otg_hpi_cs_s1_writedata                        (mm_interconnect_0_otg_hpi_cs_s1_writedata),                   //                                         .writedata
		.otg_hpi_cs_s1_chipselect                       (mm_interconnect_0_otg_hpi_cs_s1_chipselect),                  //                                         .chipselect
		.otg_hpi_data_s1_address                        (mm_interconnect_0_otg_hpi_data_s1_address),                   //                          otg_hpi_data_s1.address
		.otg_hpi_data_s1_write                          (mm_interconnect_0_otg_hpi_data_s1_write),                     //                                         .write
		.otg_hpi_data_s1_readdata                       (mm_interconnect_0_otg_hpi_data_s1_readdata),                  //                                         .readdata
		.otg_hpi_data_s1_writedata                      (mm_interconnect_0_otg_hpi_data_s1_writedata),                 //                                         .writedata
		.otg_hpi_data_s1_chipselect                     (mm_interconnect_0_otg_hpi_data_s1_chipselect),                //                                         .chipselect
		.otg_hpi_r_s1_address                           (mm_interconnect_0_otg_hpi_r_s1_address),                      //                             otg_hpi_r_s1.address
		.otg_hpi_r_s1_write                             (mm_interconnect_0_otg_hpi_r_s1_write),                        //                                         .write
		.otg_hpi_r_s1_readdata                          (mm_interconnect_0_otg_hpi_r_s1_readdata),                     //                                         .readdata
		.otg_hpi_r_s1_writedata                         (mm_interconnect_0_otg_hpi_r_s1_writedata),                    //                                         .writedata
		.otg_hpi_r_s1_chipselect                        (mm_interconnect_0_otg_hpi_r_s1_chipselect),                   //                                         .chipselect
		.otg_hpi_w_s1_address                           (mm_interconnect_0_otg_hpi_w_s1_address),                      //                             otg_hpi_w_s1.address
		.otg_hpi_w_s1_write                             (mm_interconnect_0_otg_hpi_w_s1_write),                        //                                         .write
		.otg_hpi_w_s1_readdata                          (mm_interconnect_0_otg_hpi_w_s1_readdata),                     //                                         .readdata
		.otg_hpi_w_s1_writedata                         (mm_interconnect_0_otg_hpi_w_s1_writedata),                    //                                         .writedata
		.otg_hpi_w_s1_chipselect                        (mm_interconnect_0_otg_hpi_w_s1_chipselect),                   //                                         .chipselect
		.samus_dir_s1_address                           (mm_interconnect_0_samus_dir_s1_address),                      //                             samus_dir_s1.address
		.samus_dir_s1_write                             (mm_interconnect_0_samus_dir_s1_write),                        //                                         .write
		.samus_dir_s1_readdata                          (mm_interconnect_0_samus_dir_s1_readdata),                     //                                         .readdata
		.samus_dir_s1_writedata                         (mm_interconnect_0_samus_dir_s1_writedata),                    //                                         .writedata
		.samus_dir_s1_chipselect                        (mm_interconnect_0_samus_dir_s1_chipselect),                   //                                         .chipselect
		.samus_en_s1_address                            (mm_interconnect_0_samus_en_s1_address),                       //                              samus_en_s1.address
		.samus_en_s1_write                              (mm_interconnect_0_samus_en_s1_write),                         //                                         .write
		.samus_en_s1_readdata                           (mm_interconnect_0_samus_en_s1_readdata),                      //                                         .readdata
		.samus_en_s1_writedata                          (mm_interconnect_0_samus_en_s1_writedata),                     //                                         .writedata
		.samus_en_s1_chipselect                         (mm_interconnect_0_samus_en_s1_chipselect),                    //                                         .chipselect
		.samus_jump_s1_address                          (mm_interconnect_0_samus_jump_s1_address),                     //                            samus_jump_s1.address
		.samus_jump_s1_write                            (mm_interconnect_0_samus_jump_s1_write),                       //                                         .write
		.samus_jump_s1_readdata                         (mm_interconnect_0_samus_jump_s1_readdata),                    //                                         .readdata
		.samus_jump_s1_writedata                        (mm_interconnect_0_samus_jump_s1_writedata),                   //                                         .writedata
		.samus_jump_s1_chipselect                       (mm_interconnect_0_samus_jump_s1_chipselect),                  //                                         .chipselect
		.samus_walk_s1_address                          (mm_interconnect_0_samus_walk_s1_address),                     //                            samus_walk_s1.address
		.samus_walk_s1_write                            (mm_interconnect_0_samus_walk_s1_write),                       //                                         .write
		.samus_walk_s1_readdata                         (mm_interconnect_0_samus_walk_s1_readdata),                    //                                         .readdata
		.samus_walk_s1_writedata                        (mm_interconnect_0_samus_walk_s1_writedata),                   //                                         .writedata
		.samus_walk_s1_chipselect                       (mm_interconnect_0_samus_walk_s1_chipselect),                  //                                         .chipselect
		.samus_x_s1_address                             (mm_interconnect_0_samus_x_s1_address),                        //                               samus_x_s1.address
		.samus_x_s1_write                               (mm_interconnect_0_samus_x_s1_write),                          //                                         .write
		.samus_x_s1_readdata                            (mm_interconnect_0_samus_x_s1_readdata),                       //                                         .readdata
		.samus_x_s1_writedata                           (mm_interconnect_0_samus_x_s1_writedata),                      //                                         .writedata
		.samus_x_s1_chipselect                          (mm_interconnect_0_samus_x_s1_chipselect),                     //                                         .chipselect
		.samus_y_s1_address                             (mm_interconnect_0_samus_y_s1_address),                        //                               samus_y_s1.address
		.samus_y_s1_write                               (mm_interconnect_0_samus_y_s1_write),                          //                                         .write
		.samus_y_s1_readdata                            (mm_interconnect_0_samus_y_s1_readdata),                       //                                         .readdata
		.samus_y_s1_writedata                           (mm_interconnect_0_samus_y_s1_writedata),                      //                                         .writedata
		.samus_y_s1_chipselect                          (mm_interconnect_0_samus_y_s1_chipselect),                     //                                         .chipselect
		.scene_sel_s1_address                           (mm_interconnect_0_scene_sel_s1_address),                      //                             scene_sel_s1.address
		.scene_sel_s1_write                             (mm_interconnect_0_scene_sel_s1_write),                        //                                         .write
		.scene_sel_s1_readdata                          (mm_interconnect_0_scene_sel_s1_readdata),                     //                                         .readdata
		.scene_sel_s1_writedata                         (mm_interconnect_0_scene_sel_s1_writedata),                    //                                         .writedata
		.scene_sel_s1_chipselect                        (mm_interconnect_0_scene_sel_s1_chipselect),                   //                                         .chipselect
		.sdram_s1_address                               (mm_interconnect_0_sdram_s1_address),                          //                                 sdram_s1.address
		.sdram_s1_write                                 (mm_interconnect_0_sdram_s1_write),                            //                                         .write
		.sdram_s1_read                                  (mm_interconnect_0_sdram_s1_read),                             //                                         .read
		.sdram_s1_readdata                              (mm_interconnect_0_sdram_s1_readdata),                         //                                         .readdata
		.sdram_s1_writedata                             (mm_interconnect_0_sdram_s1_writedata),                        //                                         .writedata
		.sdram_s1_byteenable                            (mm_interconnect_0_sdram_s1_byteenable),                       //                                         .byteenable
		.sdram_s1_readdatavalid                         (mm_interconnect_0_sdram_s1_readdatavalid),                    //                                         .readdatavalid
		.sdram_s1_waitrequest                           (mm_interconnect_0_sdram_s1_waitrequest),                      //                                         .waitrequest
		.sdram_s1_chipselect                            (mm_interconnect_0_sdram_s1_chipselect),                       //                                         .chipselect
		.sdram_pll_pll_slave_address                    (mm_interconnect_0_sdram_pll_pll_slave_address),               //                      sdram_pll_pll_slave.address
		.sdram_pll_pll_slave_write                      (mm_interconnect_0_sdram_pll_pll_slave_write),                 //                                         .write
		.sdram_pll_pll_slave_read                       (mm_interconnect_0_sdram_pll_pll_slave_read),                  //                                         .read
		.sdram_pll_pll_slave_readdata                   (mm_interconnect_0_sdram_pll_pll_slave_readdata),              //                                         .readdata
		.sdram_pll_pll_slave_writedata                  (mm_interconnect_0_sdram_pll_pll_slave_writedata),             //                                         .writedata
		.sysid_qsys_0_control_slave_address             (mm_interconnect_0_sysid_qsys_0_control_slave_address),        //               sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata            (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),       //                                         .readdata
		.title_en_s1_address                            (mm_interconnect_0_title_en_s1_address),                       //                              title_en_s1.address
		.title_en_s1_write                              (mm_interconnect_0_title_en_s1_write),                         //                                         .write
		.title_en_s1_readdata                           (mm_interconnect_0_title_en_s1_readdata),                      //                                         .readdata
		.title_en_s1_writedata                          (mm_interconnect_0_title_en_s1_writedata),                     //                                         .writedata
		.title_en_s1_chipselect                         (mm_interconnect_0_title_en_s1_chipselect),                    //                                         .chipselect
		.win_en_s1_address                              (mm_interconnect_0_win_en_s1_address),                         //                                win_en_s1.address
		.win_en_s1_write                                (mm_interconnect_0_win_en_s1_write),                           //                                         .write
		.win_en_s1_readdata                             (mm_interconnect_0_win_en_s1_readdata),                        //                                         .readdata
		.win_en_s1_writedata                            (mm_interconnect_0_win_en_s1_writedata),                       //                                         .writedata
		.win_en_s1_chipselect                           (mm_interconnect_0_win_en_s1_chipselect)                       //                                         .chipselect
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_qsys_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_qsys_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_qsys_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (sdram_pll_c0_clk),                       //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
