//--------------------------------------------------------------------------------------------
// Sprite Mapper:
//
//		The sprite mapper is a glorified color mapper and it will draw the sprites with the 
//		top left corner at the (x,y) coordinate. The background moves based on the position of
//		samus. (She is in the middle on the screen)
//
//--------------------------------------------------------------------------------------------
module sprite_mapper(
input logic clk, reset,
input logic vsync,
/*
// Samus
input logic enable, direction,
input logic [9:0] samus_x, samus_y,
input logic [2:0] sprite_num,

// Background
input logic scene_number,

// GUI
input logic title_en,
input logic [1:0] health,

// Monster
input logic monster1, monster2, monster3,
input logic [9:0] monster1_x, monster1_y, monster2_x, monster2_y, monster3_x, monster3_y,

// Explosion
input logic exp1_en, exp2_en, exp3_en,
input logic [9:0] exp1_x, exp1_y, exp2_x, exp2_y, exp3_x, exp3_y, 

// Bullet
input logic bullet1, bullet2, bullet3,
input logic [9:0] b1_x, b1_y, b2_x, b2_y, b3_x, b3_y,
*/

input logic [9:0] vgaX, vgaY, 
output logic [7:0] red, green, blue
);

	// Internal Signals:
	logic [6:0] bg_color;
	logic [6:0] powerUp_color;
	logic [6:0] bullet_color;
	logic [6:0] monster_color;
	logic [6:0] samus_color;
	logic [6:0] title_color;
	logic [6:0] explosion_color;
   logic [6:0] color;
	logic bulletDraw, monsterDraw, samusDraw, powerUpDraw, titleDraw, explosionDraw;
   logic [8:0] counter;
	logic [3:0] samus_temp;
 
	// This module acts as a mux on all of the different levels of sprites:
	always_ff @ (posedge vsync) begin
		counter <= counter + 1;
		if(counter >= 480) samus_temp <= 0;
		if(counter < 480) samus_temp <= 8;
		if(counter < 450) samus_temp <= 15;
		if(counter < 420) samus_temp <= 7;
		if(counter < 390) samus_temp <= 14;
		if(counter < 360) samus_temp <= 6;
		if(counter < 330) samus_temp <= 13;
		if(counter < 300) samus_temp <= 5;
		if(counter < 270) samus_temp <= 12;
		if(counter < 240) samus_temp <= 4;
		if(counter < 210) samus_temp <= 11;
		if(counter < 180) samus_temp <= 3;
		if(counter < 150) samus_temp <= 10;
		if(counter < 120) samus_temp <= 2;
		if(counter < 90) samus_temp <= 9;
		if(counter < 60) samus_temp <= 1;
		if(counter < 30) samus_temp <= 1;
	end
	
	
	
   // Texture Units: 
	
	background bg(.background_start_addr(1'b0), .vga_x(vgaX), .vga_y(vgaY), .color(bg_color)); 
   bullet bull(.enable1(1'b1), .enable2(1'b1), .enable3(1'b1), 
		.vga_x(vgaX), .vga_y(vgaY), 
		.sprite1_x(120), .sprite1_y(40), 
		.sprite2_x(80), .sprite2_y(40), 
		.sprite3_x(40), .sprite3_y(40), 
		.empowered(1'b1),
		.color(bullet_color),
		.draw(bulletDraw));
	monster mon(.enable1(1'b1), .enable2(1'b1), .enable3(1'b1),
					.vga_x(vgaX), .vga_y(vgaY), 
					.sprite1_x(40), .sprite1_y(80), 
					.sprite2_x(100), .sprite2_y(80), 
					.sprite3_x(160), .sprite3_y(80),
					.color(monster_color), .draw(monsterDraw)); 
	samus(.enable(1'b1), .vga_x(vgaX), .vga_y(vgaY),
			.sprite_x(40), .sprite_y(140), .sprite_num(samus_temp[2:0]),
			.direction(samus_temp[3]), .color(samus_color), .draw(samusDraw));
	gui info(.titleEn(1'b0), .health(samus_temp[1:0]),
				.vga_x(vgaX), .vga_y(vgaY),
				.color(title_color), .draw(titleDraw));
	explosion explode(.enable1(samus_temp[0]), .enable2(samus_temp[1]), .enable3(samus_temp[2]), .vsync(vsync), 
							.vga_x(vgaX), .vga_y(vgaY), 
							.exp1_x(240), .exp1_y(40), 
							.exp2_x(340), .exp2_y(40), 
							.exp3_x(440), .exp3_y(40),
							.color(explosion_color), .draw(explosionDraw));
	
	
	// Select the color based on priority:
	always_comb begin
	   // Default:
	   color = bg_color;
	   if(titleDraw == 1'b1) color = title_color;
		else if(explosionDraw == 1'b1) color = explosion_color;
		else if(samusDraw == 1'b1) color = samus_color;
		else if(monsterDraw == 1'b1) color = monster_color;
		else if(bulletDraw == 1'b1) color = bullet_color;
		else color = bg_color; 
	end
	
	// Pass the color to pallate to output the proper color:
	always_comb begin
		//Defaults:
		red = 8'b0;
		green = 8'b0;
		blue = 8'b0;
		
		case(color)
			//Color 1:
			1: begin
				red = 44;
				green = 92;
				blue = 10;
			end
			//Color 2:
			2: begin
			//248,146,56
				red = 248;
				green = 146;
				blue = 56;
			end
			//Color 3:
			3: begin
			//(156,0,18
				red = 156;
				green = 0;
				blue = 18;
			end
			//Color 4:
			4: begin
			// 0, 255, 128
				red = 0;
				green = 255;
				blue = 128;
			end
			//Color 5:
			5: begin
			// 0,0,128
				red = 0;
				green = 0;
				blue = 128;
			end
			//Color 6:
			6: begin
			// 0,128,255
				red = 0;
				green = 128;
				blue = 255;
			end
			//Color 7:
			7: begin
			// 255,255,255
				red = 255;
				green = 255;
				blue = 255;
			end
			//Color 8:
			8: begin
				red = 0;
				green = 0;
				blue = 0;
			end
			//Color 9:
			9: begin
				red = 0;
				green = 0;
				blue = 255;
			end
			//Color 10:
			10: begin
				red = 102;
				green = 102;
				blue = 102;
			end
			//Color 11:
			11: begin
				red = 0;
				green = 255;
				blue = 255;
			end
			//Color 12
			12: begin
				red = 0;
				green = 255;
				blue = 0;
			end
			//Color 13:
			13: begin
				red = 64;
				green = 128;
				blue = 0;
			end
			//Color 14:
			14: begin
				red = 255;
				green = 0;
				blue = 0;
			end
			//Color 15:
			15: begin
				red = 255;
				green = 102;
				blue = 102;
			end
			//Color 16
			16: begin
				red = 128;
				green = 0;
				blue = 0;
			end
			//Color 17:
			17: begin
				red = 248;
				green = 146;
				blue = 56;
			end
			//Color 18:
			18: begin
				red = 232;
				green = 146;
				blue = 41;
			end
			//Color 19:
			19: begin
				red = 27;
				green = 175;
				blue = 0;
			end
			//Color 20:
			20: begin
				red = 19;
				green = 137;
				blue = 13;
			end
			//Color 21:
			21: begin
				red = 255;
				green = 49;
				blue = 62;
			end
			//Color 22:
			22: begin
				red = 234;
				green = 228;
				blue = 94;
			end
			//Color 23:
			23: begin
				red = 126;
				green = 0;
				blue = 246;
			end
			//Color 24:
			24: begin
				red = 47;
				green = 151;
				blue = 209;
			end
			//Color 25:
			25: begin
				red = 156;
				green = 89;
				blue = 33;
			end
			//Color 26:
			26: begin
				red = 82;
				green = 105;
				blue = 250;
			end
			//Color 27:
			27: begin
				red = 43;
				green = 93;
				blue = 83;
			end
			//Color 28:
			28: begin
				red = 13;
				green = 65;
				blue = 63;
			end
			//Color 29:
			29: begin
				red = 37;
				green = 75;
				blue = 258;
			end
			//Color 30:
			30: begin
				red = 148;
				green = 148;
				blue = 118;
			end
			//Color 31:
			31: begin
				red = 60;
				green = 70;
				blue = 17;
			end
			//Color 32:
			32: begin
				red = 63;
				green = 71;
				blue = 73;
			end
			//Color 33:
			33: begin
				red = 34;
				green = 28;
				blue = 28;
			end
			34: begin
				red = 4;
				green = 35;
				blue = 248;
			end
			35: begin
				red = 186;
				green = 0;
				blue = 37;
			end
			36: begin
				red = 103;
				green = 0;
				blue = 246;
			end
			37: begin
				red = 103;
				green = 0;
				blue = 183;
			end
			// Default:
			default: begin
				red = 0;
				green = 0;
				blue = 0;
			end
		endcase
	end
	
endmodule



//--------------------------------------------------------------------------------------------
// Samus:
//
//		If the vga pixel pointer is within the samus sprite, return a proper color:
//		Priority 1
//
//--------------------------------------------------------------------------------------------
module samus(
	input logic  			enable,
	input logic  [10:0] 	vga_x, vga_y, sprite_x, sprite_y,
	input logic  [2:0] 	sprite_num,
	input logic direction,
	output logic [5:0] 	color,
	output logic 			draw
);
   // Direction:
   // 0 is right
	// 1 is left

	// Samus Sprites:
	parameter [9:0] height1 = 69;
	parameter [9:0] width1 = 45;
	
	parameter [9:0] height2 = 69;
	parameter [9:0] width2 = 45;
	
	parameter [9:0] height3 = 70;
	parameter [9:0] width3 = 45;
	
	parameter [9:0] height4 = 58;
	parameter [9:0] width4 = 45;
	
	parameter [9:0] height5 = 57;
	parameter [9:0] width5 = 45;
	
	parameter [9:0] height6 = 54;
	parameter [9:0] width6 = 45;
	
	parameter [9:0] height7 = 68;
	parameter [9:0] width7 = 45;
	
	// Sprites:
	int samus1[height1][width1];
	int samus2[height2][width2];
	int samus3[height3][width3];
	int samus4[height4][width4];
	int samus5[height5][width5];
	int samus6[height6][width6];
	int samus7[height7][width7];
	
	always_ff begin
		// Samus Standing Up:
		samus1 =  '{'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,31,31,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,31,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,31,31,31,19,31,1,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,31,25,31,31,19,31,25,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,18,31,1,25,25,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,25,25,31,19,31,25,25,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,31,19,31,31,31,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,31,31,31,19,31,19,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,31,19,31,31,31,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,18,18,25,25,1,25,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,2,18,31,25,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,3,3,3,18,2,18,2,2,18,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,33,33,33,16,3,3,3,18,2,2,2,2,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,3,35,3,3,3,21,3,18,2,2,2,18,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,33,16,3,3,3,21,3,3,3,21,21,18,18,21,21,21,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,3,3,3,21,3,3,3,3,3,3,3,2,21,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,16,3,3,3,3,3,21,31,31,18,18,21,3,3,3,3,3,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,3,3,21,3,3,3,3,25,31,18,18,3,3,21,3,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,16,3,18,2,3,3,21,31,25,1,31,18,2,2,21,3,21,18,21,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,16,3,18,2,3,3,21,31,31,25,25,18,2,2,18,21,21,18,21,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,16,3,18,2,3,21,18,25,31,25,2,2,2,2,18,2,25,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,16,3,21,21,3,21,18,25,25,25,2,2,2,2,2,2,21,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,16,3,3,3,3,21,18,25,31,18,2,2,2,2,2,18,21,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,33,3,3,18,21,2,25,31,18,18,2,2,18,18,25,25,3,16,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,3,3,18,2,2,25,31,18,2,2,2,2,18,31,31,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,2,2,2,18,18,2,2,2,2,2,21,16,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,18,2,2,2,2,2,2,2,18,2,18,3,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,18,2,2,2,2,2,2,2,18,31,31,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,2,2,2,2,2,2,2,2,18,31,31,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,18,2,2,2,18,2,18,2,18,31,31,3,21,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,31,31,2,2,2,2,2,2,18,31,31,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,33,2,18,2,2,2,18,2,31,31,3,21,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,33,2,2,2,2,2,2,2,18,25,31,16,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,33,2,2,2,2,2,2,2,18,18,31,25,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,33,2,18,2,2,2,18,2,2,2,18,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,18,2,18,2,2,2,2,2,2,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,31,2,2,2,2,2,2,18,2,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,2,2,2,18,2,2,18,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,31,2,2,2,2,2,2,25,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,25,25,2,2,18,2,2,18,25,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,33,18,2,2,2,2,2,2,2,25,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,33,2,2,2,2,2,2,2,2,18,18,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,33,2,2,2,2,2,2,2,2,2,2,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,33,2,2,2,2,2,2,2,2,18,2,2,18,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,25,18,2,2,2,2,2,2,2,2,2,2,31,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,31,2,2,18,2,2,18,2,2,2,2,2,18,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,2,2,2,2,18,31,25,18,2,2,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,31,2,2,2,2,18,33,33,2,2,18,2,18,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,31,18,2,18,2,18,33,33,33,25,2,21,16,3,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,31,2,2,2,2,18,33,33,33,31,2,21,3,3,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,2,2,2,2,18,33,33,33,31,2,2,2,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,31,2,2,18,18,21,33,33,33,25,2,2,2,16,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,31,18,2,2,3,3,3,21,18,2,2,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,25,2,21,21,3,3,3,21,18,2,2,25,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,33,2,2,2,21,3,21,3,3,21,18,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,25,25,2,2,2,18,21,16,21,21,18,2,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,2,2,2,2,2,2,2,3,3,18,2,18,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,16,3,25,18,2,2,18,2,2,31,0,33,33,2,2,2,21,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,16,3,18,2,18,18,18,18,18,16,0,0,33,18,2,18,21,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,33,3,3,3,18,18,3,3,3,16,0,0,0,3,3,2,21,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,33,3,3,3,21,21,3,3,16,16,0,0,0,3,3,18,21,3,16,25,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,33,35,3,21,3,3,21,16,0,0,0,0,0,3,3,3,3,3,25,31,16,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,33,3,3,3,25,31,31,31,0,0,0,0,0,3,3,3,25,31,31,31,3,3,16,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,33,3,21,3,31,31,31,31,0,0,0,0,0,3,3,3,16,25,31,3,21,3,3,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,33,33,31,16,16,25,16,3,33,0,0,0,0,33,3,25,31,25,3,3,3,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,33,25,16,3,3,3,3,16,0,0,0,0,0,3,16,31,31,3,3,21,3,3,3,16,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}};
		
		// Running Forward 1:
		samus2 =  '{'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,16,16,16,16,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,3,3,3,3,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,3,3,3,3,21,3,3,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,3,3,21,3,3,3,3,3,3,3,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,18,2,3,3,3,3,3,21,3,3,21,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,33,3,21,21,21,3,3,21,16,25,3,3,3,16,25,21,25,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,16,3,2,18,3,3,3,3,3,31,31,3,21,3,25,31,25,18,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,16,3,21,21,3,3,21,3,3,25,31,25,31,3,16,33,31,25,31,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,16,3,3,3,3,3,3,3,21,3,3,31,31,3,16,33,31,31,18,18,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,16,3,3,21,3,21,3,3,3,25,31,16,16,3,16,33,31,1,25,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,16,3,3,3,3,3,3,21,3,31,31,3,21,3,16,33,31,31,31,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,18,18,2,18,2,31,33,16,3,3,3,3,3,3,33,33,1,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,18,18,2,31,33,16,3,3,3,21,3,3,16,33,31,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,33,31,18,2,31,25,2,2,2,33,33,3,3,3,3,3,3,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,31,25,2,18,25,18,18,2,2,31,31,21,21,21,21,3,21,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,25,2,2,2,2,2,2,2,2,2,2,18,2,18,21,3,3,3,21,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,33,25,18,2,25,25,2,2,2,18,2,18,2,25,31,31,31,31,16,3,21,18,25,25,25,31,31,31,33,25,31,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,31,18,2,2,31,31,2,2,2,2,2,2,2,31,1,33,33,25,16,21,18,18,18,18,2,25,1,31,31,18,18,31,31,0,0,0},
						'{0,0,0,0,0,0,0,0,0,31,2,2,2,25,31,18,2,2,2,2,2,2,18,18,18,18,18,18,18,18,2,2,2,2,25,31,19,31,25,31,1,31,1,0,0},
						'{0,0,0,0,0,0,0,0,0,16,18,18,2,31,25,2,2,18,2,18,2,2,2,2,2,2,2,18,18,2,2,2,2,18,25,31,31,1,25,1,25,1,25,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,25,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,21,3,18,2,2,18,31,31,19,31,25,1,25,1,25,1,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,31,25,25,25,2,2,2,2,2,2,2,18,2,2,18,2,21,3,21,21,25,31,25,1,31,31,19,25,25,1,31,1,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,18,2,2,2,2,2,2,2,2,18,25,3,3,16,33,33,31,25,1,25,1,2,18,31,31,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,2,2,2,2,2,18,2,2,2,2,21,21,3,3,25,31,33,33,33,33,33,31,31,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,2,2,2,2,2,2,2,2,2,2,2,2,21,3,18,25,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,2,2,2,2,2,2,18,33,25,18,2,2,3,21,2,25,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,2,2,2,2,2,18,18,33,31,2,2,2,3,16,2,25,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,2,2,2,2,2,2,25,33,33,33,16,3,2,18,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,2,2,2,2,2,2,2,2,18,33,33,33,16,21,18,21,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,18,2,2,2,18,2,2,18,2,18,2,2,21,21,21,25,16,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,2,2,2,2,2,2,2,2,2,2,2,2,21,3,18,2,2,25,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,2,2,2,2,2,2,18,2,2,2,25,16,25,21,2,2,2,25,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,18,18,2,2,2,2,2,2,2,2,18,2,31,33,25,2,2,2,18,25,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,2,2,2,2,18,0,33,33,33,33,31,18,18,2,2,18,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,2,2,2,33,33,33,33,33,31,2,18,18,18,18,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,2,18,2,33,33,3,3,2,2,2,21,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,2,18,25,16,33,3,21,21,21,18,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,2,31,0,16,3,3,3,3,3,3,21,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,31,25,18,2,2,31,0,3,3,3,21,31,25,31,16,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,18,18,2,2,2,31,0,16,3,3,16,25,1,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,33,25,25,18,21,16,2,25,33,0,0,3,3,25,31,16,16,25,3,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,31,2,2,18,3,21,2,25,0,0,0,16,3,31,31,3,3,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,16,3,3,3,2,2,2,2,2,3,3,3,16,0,0,0,0,0,0,33,3,21,3,3,21,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,3,3,3,21,2,2,18,2,2,21,3,16,16,0,0,0,0,0,0,0,3,3,3,3,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,16,3,3,3,3,21,18,2,2,2,18,3,3,0,0,0,0,0,0,0,0,0,0,33,3,21,3,3,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,33,25,31,25,3,3,21,21,21,25,31,16,16,0,0,0,0,0,0,0,0,0,0,33,16,16,16,16,16,16,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,33,31,31,31,3,21,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,33,31,16,25,31,31,3,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,16,3,3,3,25,31,3,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,16,3,21,3,3,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,16,3,3,3,3,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,16,3,3,21,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,16,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,16,3,21,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,16,16,3,3,3,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,3,3,3,3,3,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,33,33,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}};
		
		// Running Forward 2:
		samus3 =  '{'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,3,3,3,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,3,3,3,3,3,3,3,3,3,3,3,3,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,16,21,3,3,3,21,3,21,3,3,3,3,3,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,3,21,18,21,3,3,3,3,3,3,21,3,21,3,3,3,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,16,21,21,25,3,21,3,21,31,25,3,3,3,31,25,21,16,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,21,18,21,3,3,3,3,16,31,31,3,21,3,31,31,2,25,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,25,3,3,3,21,3,3,25,16,31,16,3,33,33,25,31,18,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,3,3,21,3,3,3,3,3,25,31,25,3,33,33,31,25,2,31,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,21,3,3,3,3,21,16,25,31,3,3,3,33,33,1,31,31,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,3,3,3,21,3,3,16,31,31,3,3,3,33,33,31,1,25,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,3,3,3,3,3,21,3,3,3,21,3,3,3,3,33,33,1,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,21,21,21,21,21,25,21,16,3,3,3,21,3,3,16,16,31,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,18,2,2,18,18,18,25,33,16,3,3,3,3,3,3,3,3,16,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,33,25,25,25,25,25,25,25,2,25,25,18,2,2,18,33,33,3,3,21,3,3,16,33,16,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,31,18,18,18,18,2,18,2,2,25,31,18,2,2,25,33,16,3,3,3,3,3,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,3,3,3,25,25,33,33,33,31,2,2,18,2,2,2,21,3,16,33,16,3,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,3,21,16,25,31,33,33,33,16,18,18,18,18,18,18,18,16,16,33,3,21,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,33,2,2,2,2,2,2,2,2,25,25,1,25,1,25,1,25,31,25,2,18,2,18,18,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,33,2,2,2,2,2,2,2,2,18,25,25,1,25,1,31,31,1,25,18,18,2,2,18,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,33,2,2,2,2,2,2,18,2,2,18,25,31,31,19,31,19,31,31,25,25,2,2,2,2,25,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,31,25,2,2,2,2,2,2,2,2,25,1,31,33,33,33,33,1,1,18,2,18,2,2,25,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,31,2,2,2,2,2,2,2,2,25,25,33,33,33,33,33,33,31,18,18,2,2,18,25,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,33,33,33,18,2,2,18,25,31,1,1,31,31,31,31,31,18,18,2,2,18,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,2,18,31,19,31,25,1,31,31,19,25,2,2,2,2,18,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,2,2,2,2,2,18,18,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,2,2,18,2,2,18,18,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,2,2,2,2,2,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,25,2,2,18,2,2,21,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,2,2,2,2,18,2,18,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,16,16,16,16,16,33,0,0,0,0,0,2,2,2,18,2,2,2,2,25,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,16,3,3,3,3,16,0,0,0,0,0,18,2,2,2,2,2,18,2,18,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,33,1,16,21,3,3,21,16,0,0,0,0,0,18,2,2,18,2,2,2,2,18,18,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,33,31,16,3,3,3,3,16,0,0,0,0,0,18,18,2,2,2,2,18,2,2,2,25,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,33,3,3,3,31,25,3,21,3,3,3,33,0,0,0,0,33,2,2,2,2,2,2,2,18,18,18,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,33,3,3,21,31,31,3,3,21,21,21,16,33,0,0,33,25,18,2,2,25,25,2,2,2,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,33,35,3,3,31,31,16,21,18,18,18,2,2,0,0,18,2,2,2,2,33,0,18,2,2,2,2,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,16,16,3,3,3,31,33,3,21,25,21,2,2,2,16,16,2,2,18,25,31,0,0,31,31,2,18,2,25,31,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,3,3,21,3,3,33,0,3,3,3,21,2,2,18,3,21,18,2,2,31,0,0,0,0,33,2,2,2,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,3,3,3,16,33,0,0,33,16,3,21,18,2,2,3,21,18,2,2,31,0,0,0,0,33,2,2,2,2,18,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,3,3,3,16,0,0,0,0,0,3,21,18,2,2,3,16,18,2,2,31,0,0,0,0,33,2,18,2,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,25,2,18,2,3,3,0,0,0,0,0,0,0,0,16,3,3,3,3,3,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,31,18,18,21,3,16,0,0,0,0,0,0,0,0,33,21,21,21,3,3,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,3,16,0,0,0,0,0,0,0,0,16,18,18,18,3,3,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,16,16,33,0,0,0,0,0,0,0,31,25,2,2,2,16,16,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,18,2,2,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,25,25,2,2,2,31,16,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,2,2,2,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,3,2,2,18,21,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,18,18,18,21,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,3,3,3,3,3,3,3,3,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,3,3,3,21,3,25,16,25,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,3,21,3,3,16,25,31,31,31,3,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,16,3,25,31,31,31,25,3,3,16,16,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,31,31,3,3,3,3,3,3,3,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,0,33,3,21,3,21,3,3,3,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,3,3,3,3,3,21,3,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}};
		
		// Running Forward 3:
		samus4 =  '{'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,3,3,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,33,33,16,3,3,3,3,3,33,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,35,3,3,21,3,3,3,3,3,3,35,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,16,21,21,3,3,3,3,21,3,3,21,3,3,3,16,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,16,2,21,3,3,21,3,3,3,3,3,3,3,3,3,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,16,21,18,21,16,3,3,3,25,31,3,21,3,25,31,18,18,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,3,2,18,3,3,21,3,3,31,25,3,3,3,25,31,18,18,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,3,3,3,3,3,3,3,21,3,3,25,31,3,16,33,31,31,18,18,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,3,21,3,16,3,16,3,3,16,16,31,31,3,16,33,31,1,18,18,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,3,3,3,33,33,33,16,3,31,25,3,3,21,16,33,31,31,31,1,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,16,3,3,31,31,31,25,21,31,31,3,3,3,16,16,33,33,1,31,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,21,18,2,18,18,2,33,33,3,3,3,3,3,33,33,1,1,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,31,31,2,18,25,18,2,25,25,33,16,3,3,3,16,16,16,16,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,31,2,18,31,25,2,2,2,33,33,3,21,3,3,3,3,3,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,2,18,18,25,25,18,2,31,31,3,3,3,21,3,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,2,2,2,25,31,18,18,31,31,3,21,3,3,3,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,25,18,2,2,2,2,2,2,2,25,31,3,25,31,31,3,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,18,18,2,18,25,25,25,25,25,25,25,21,16,31,31,16,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,31,2,2,2,2,18,33,33,33,33,33,25,2,2,18,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,21,21,21,18,18,31,31,31,31,31,21,21,25,21,16,33,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,3,3,3,2,2,2,2,2,2,2,3,3,3,3,3,31,31,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,3,21,18,18,2,2,2,2,21,21,3,3,31,31,31,31,25,1,31,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,3,21,2,2,2,2,2,2,21,3,3,21,31,31,25,1,31,31,31,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,25,2,2,2,18,2,18,21,3,33,33,33,33,33,33,33,1,1,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,31,18,18,2,2,2,2,21,16,16,33,33,33,33,33,33,33,1,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,2,2,2,2,2,3,3,3,3,31,31,31,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,18,2,2,2,2,16,16,16,16,31,28,31,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,2,2,18,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,25,18,2,2,2,2,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,25,18,2,2,18,2,2,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,25,2,2,2,2,2,18,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,25,18,2,2,2,2,2,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,25,18,2,2,18,2,2,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,31,25,18,2,2,2,2,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,2,18,2,21,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,2,2,2,21,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,18,2,2,21,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,2,2,18,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,2,2,2,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,3,3,3,3,3,2,21,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,33,16,3,21,3,21,21,18,18,21,16,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,3,3,3,3,3,21,18,2,18,2,2,18,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,33,16,3,3,25,25,21,18,2,2,2,2,18,25,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,16,3,3,25,31,25,18,2,2,2,2,2,25,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,3,3,3,21,25,18,2,2,18,2,18,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,16,3,3,21,18,2,2,2,2,2,18,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,18,18,2,2,2,21,3,3,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}};
		
		// Jumping Up:
		samus5 =  '{'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,31,1,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,31,31,25,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,31,19,31,1,31,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,25,25,31,31,19,25,25,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,18,31,19,31,18,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,25,25,31,31,31,25,25,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,31,19,31,1,25,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,31,31,31,19,31,31,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,25,1,31,25,1,25,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,18,25,31,19,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,18,2,2,18,25,31,25,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,3,3,35,18,2,2,2,2,2,18,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,16,33,3,3,3,3,2,2,2,18,2,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,3,3,3,21,3,18,2,2,2,2,2,18,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,16,16,3,3,3,21,3,3,3,21,21,18,21,21,21,21,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,3,21,3,3,3,3,3,3,21,18,21,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,3,3,3,3,21,31,31,2,21,16,3,3,3,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,3,21,3,3,21,3,3,31,25,2,18,21,3,21,3,21,3,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,16,3,18,18,3,3,3,25,31,31,1,18,2,18,21,3,18,18,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,16,3,18,18,3,21,21,31,19,25,25,2,2,2,21,21,21,21,16,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,16,3,2,18,3,21,18,25,31,18,2,2,2,2,2,18,25,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,16,3,21,21,3,21,18,25,31,18,2,2,2,2,2,18,21,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,16,3,3,3,3,21,18,25,31,18,2,18,2,2,2,2,21,3,21,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,33,3,21,18,18,2,25,31,18,2,2,2,18,18,25,16,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,2,2,2,25,31,18,2,2,2,2,25,31,25,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,2,2,18,2,2,18,2,2,21,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,2,2,2,2,2,2,2,18,25,3,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,2,18,2,2,18,2,18,1,25,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,2,2,2,2,2,2,18,31,31,3,21,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,2,2,18,2,2,18,18,31,31,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,31,2,2,2,2,2,2,18,31,31,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,2,2,18,2,2,2,18,31,25,3,21,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,2,2,2,2,2,2,2,18,25,31,16,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,2,2,2,2,2,2,2,2,25,25,31,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,2,2,18,2,2,2,18,2,2,2,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,25,18,2,2,18,2,2,2,2,2,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,31,2,2,2,2,2,2,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,31,2,2,2,2,18,2,25,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,31,2,2,2,2,2,2,25,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,16,16,3,16,0,33,25,18,2,2,18,2,2,18,18,25,25,25,25,25,25,25,16,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,16,3,3,3,0,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,21,3,16,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,3,16,31,31,3,3,3,0,33,2,2,2,2,2,2,2,2,2,2,2,2,2,18,3,21,2,2,18,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,16,3,31,31,25,16,21,3,0,16,25,2,2,2,2,2,2,2,2,2,18,2,18,18,21,25,18,2,2,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,3,3,3,3,3,25,31,16,3,3,16,33,31,2,2,2,18,2,2,18,2,2,2,33,33,18,18,2,2,2,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,3,3,21,3,3,31,31,16,21,21,16,33,31,2,2,2,2,18,31,25,31,25,31,31,31,2,2,2,25,25,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,3,3,3,3,21,31,25,3,3,18,25,33,31,2,2,2,18,18,33,33,33,33,33,18,2,2,2,2,31,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,3,3,16,33,33,16,16,3,21,2,18,25,25,21,18,18,2,25,33,33,16,31,25,18,18,21,16,31,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,3,16,0,0,0,16,3,3,21,18,2,2,21,3,18,2,2,18,33,16,3,21,2,2,18,3,16,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,18,2,2,21,3,21,2,0,33,3,3,3,3,21,3,21,3,16,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,16,3,2,18,2,21,3,18,2,0,0,3,3,3,21,16,3,16,3,16,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,2,2,2,2,2,0,33,3,3,3,31,31,25,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,21,21,21,25,25,0,0,3,21,31,25,31,31,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,3,3,3,33,0,0,33,3,31,31,16,3,3,3,3,16,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,16,16,0,0,0,0,16,33,31,16,3,21,3,3,3,16,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,3,3,3,21,3,3,16,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,3,3,3,3,3,3,16,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,21,3,3,3,3,0,0,0,0,0,0,0,0,0}};
		
		// Jumping Moving:
		samus6 =  '{'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,3,3,35,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,33,16,3,3,3,3,3,16,16,33,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,3,3,3,3,3,21,3,3,3,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,16,21,21,3,3,3,3,3,21,3,3,3,3,16,16,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,35,21,2,21,3,21,3,21,3,3,3,21,3,3,3,16,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,2,21,3,3,3,3,16,31,31,3,3,3,25,25,18,25,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,21,18,21,3,3,21,3,3,25,31,21,3,3,31,1,2,25,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,3,3,3,3,3,3,3,3,25,1,25,3,33,33,31,25,18,31,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,3,3,16,16,16,3,21,16,31,31,16,3,33,33,1,25,18,31,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,21,16,33,33,33,3,16,25,31,3,21,3,33,33,31,31,31,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,16,3,16,31,31,31,21,25,33,31,3,3,3,16,16,33,31,1,31,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,21,2,2,2,2,18,33,33,3,3,3,3,3,33,33,31,31,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,25,18,21,18,2,2,2,18,18,18,21,18,18,18,21,3,16,16,18,31,31,31,31,25,25,31,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,21,2,25,31,31,1,18,2,1,31,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,25,2,2,2,2,2,2,2,2,2,18,31,25,2,2,2,18,2,18,2,2,25,25,1,25,31,31,19,31,1,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,21,2,2,2,2,2,2,2,18,18,18,25,25,2,2,2,2,2,2,2,18,25,31,19,31,1,25,1,25,31,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,16,3,18,2,2,2,2,2,2,2,2,31,31,2,2,2,2,2,2,2,2,18,31,31,31,31,19,31,31,31,1,25,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,16,3,18,18,2,2,18,2,2,18,25,25,25,18,2,21,18,2,2,2,2,18,1,33,1,1,31,25,25,25,1,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,16,3,2,2,2,2,2,2,2,25,31,18,2,2,21,3,21,2,18,2,2,25,0,0,0,31,31,18,18,31,1,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,33,21,2,2,18,2,2,2,18,25,2,2,25,25,3,21,21,16,31,16,33,0,0,0,0,33,33,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,25,2,2,2,2,2,2,2,2,2,18,31,31,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,2,2,2,2,2,2,2,18,18,31,31,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,18,2,2,2,2,2,2,2,2,18,31,25,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,2,2,2,2,2,2,2,18,2,2,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,2,2,2,2,2,2,2,2,18,25,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,2,2,2,2,2,18,2,2,25,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,16,16,16,0,0,31,25,18,2,2,18,2,2,2,18,18,31,31,31,31,31,16,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,33,3,3,3,0,0,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,16,16,31,31,3,3,3,33,0,2,2,2,2,2,2,2,2,2,2,2,2,2,2,21,3,18,18,25,31,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,3,3,31,31,3,21,3,33,0,18,2,2,2,2,2,2,2,18,2,2,18,2,18,21,3,18,2,2,31,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,16,3,3,3,3,25,31,31,3,3,3,33,33,2,2,2,2,2,2,2,2,2,2,31,33,25,2,2,2,2,31,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,3,3,3,21,3,16,25,31,3,21,3,33,33,2,2,18,2,2,18,25,18,18,25,31,33,18,2,2,18,18,31,0,0,0,0,0,0,0,0,0,0},
						'{0,0,16,3,3,3,3,3,3,25,31,31,3,18,18,33,33,2,2,2,2,2,33,33,33,33,33,31,2,2,2,2,18,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,33,3,3,21,16,16,16,16,31,16,3,18,2,31,31,21,21,2,2,18,33,33,33,16,31,18,2,21,21,31,31,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,16,3,3,3,0,0,0,33,3,3,21,21,2,2,21,3,21,2,2,2,33,33,3,21,18,18,2,21,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,33,16,33,0,0,0,0,16,16,3,18,2,2,18,3,21,18,31,16,16,3,3,3,21,21,16,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,16,3,18,18,2,18,3,21,2,16,0,3,3,3,3,3,3,3,21,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,18,2,18,18,2,33,0,3,3,21,16,25,31,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,18,18,18,18,18,16,0,3,3,16,25,31,31,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,3,16,0,0,0,3,16,25,31,3,3,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,16,3,33,0,0,0,16,16,31,31,3,3,21,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,3,3,3,3,21,3,3,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,16,3,3,3,3,3,16,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,16,3,21,3,3,3,3,16,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,0,33,33,0,0,0,0,0,0,0,0,0,0,0,0,0}};
						
		samus7 =  '{'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,33,33,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,35,3,35,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,33,16,16,16,3,3,3,3,3,16,16,16,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,16,3,3,3,3,3,21,3,3,3,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,16,25,21,21,3,3,3,3,3,21,3,3,21,3,16,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,35,21,18,21,3,21,3,21,3,3,3,3,3,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,3,21,18,21,3,3,3,3,16,31,31,3,21,3,31,25,2,18,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,3,3,18,21,3,3,21,3,3,31,25,16,3,3,31,31,18,25,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,3,3,3,3,3,3,3,3,21,3,31,25,31,3,33,33,31,25,18,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,3,3,21,3,3,21,3,3,3,25,16,31,16,3,33,33,1,31,18,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,3,3,3,3,3,3,3,21,3,31,31,3,21,3,33,33,31,31,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,33,16,3,21,21,18,21,21,18,18,25,33,16,3,3,16,33,33,19,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,33,3,21,2,2,2,2,2,2,25,33,16,3,3,3,33,33,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,33,18,18,2,2,2,2,18,31,25,18,31,33,3,3,3,16,16,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,33,2,2,2,2,2,18,18,31,25,18,31,33,16,3,21,3,21,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,18,2,2,2,2,18,2,31,25,18,25,31,25,2,21,3,18,2,2,2,2,31,31,1,31,2,18,1,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,18,2,2,2,2,18,18,25,25,18,18,25,18,18,21,21,2,2,2,2,2,25,31,25,31,25,25,31,31,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,18,2,2,18,2,25,1,2,2,2,2,2,2,2,18,18,18,2,2,18,2,25,31,1,25,31,19,31,31,1,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,18,2,2,2,2,31,33,18,2,2,2,18,21,21,21,25,18,2,2,18,25,31,19,31,1,25,1,25,1,25,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,18,2,2,2,2,16,33,18,2,2,2,2,21,3,3,3,2,2,2,25,31,25,1,25,31,1,25,1,25,1,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,18,2,2,2,2,18,25,25,25,16,21,18,18,18,21,3,21,16,33,31,31,1,25,1,25,18,25,31,1,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,18,2,2,18,2,2,2,31,31,3,21,18,2,18,3,3,3,16,0,33,19,31,31,31,25,18,18,1,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,33,2,2,2,2,2,25,31,3,3,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,33,2,2,18,2,2,25,31,3,21,3,21,21,33,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,33,2,2,2,2,18,2,18,3,3,3,21,18,3,3,3,35,3,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,31,18,18,2,2,2,18,25,25,31,18,2,21,21,3,3,3,16,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,31,2,2,2,2,18,31,31,31,25,2,2,2,3,21,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,16,2,2,18,2,2,18,31,33,33,16,16,21,3,3,33,16,3,16,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,31,2,2,2,2,2,2,25,0,0,0,3,3,3,16,0,16,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,18,18,2,2,2,18,2,2,25,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,33,2,2,18,2,2,2,2,18,25,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,33,2,2,2,2,2,2,2,2,2,18,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,33,2,2,2,2,2,2,2,2,2,2,25,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,33,2,2,2,2,2,2,2,18,2,18,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,31,25,2,2,2,2,2,2,2,2,2,2,25,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,31,2,2,2,2,2,2,2,2,18,2,18,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,31,2,2,2,2,18,33,31,2,2,2,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,16,2,2,18,2,18,33,16,2,2,2,18,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,31,2,2,2,2,18,33,33,33,31,2,21,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,31,18,2,2,2,18,33,33,33,31,2,21,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,31,2,2,18,2,18,33,33,33,31,2,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,16,2,2,2,21,21,33,16,31,25,2,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,31,2,2,2,3,3,3,21,18,2,2,2,18,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,25,25,2,21,21,3,3,3,21,18,2,2,31,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,0,33,18,2,2,21,3,3,21,3,21,18,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,18,18,2,2,2,18,18,3,21,18,18,2,18,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,0,0,0,0,18,2,2,2,2,18,18,16,16,2,2,2,18,18,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,16,3,21,2,2,2,18,2,2,16,0,0,0,2,2,2,21,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,33,16,3,18,2,21,21,21,18,25,33,0,33,16,2,18,21,21,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,33,3,3,3,18,2,3,3,3,16,0,0,0,3,3,2,21,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,33,35,3,21,21,25,3,3,16,0,0,0,0,3,3,21,21,3,25,31,16,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,33,3,3,3,3,3,3,16,0,0,0,0,0,3,3,3,16,3,31,31,16,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,33,3,3,3,25,31,31,31,0,0,0,0,0,3,3,3,25,31,25,16,3,3,3,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,33,3,21,3,31,31,31,1,0,0,0,0,0,3,3,3,16,25,16,3,21,3,3,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,33,31,16,3,3,3,3,16,0,0,0,0,0,3,25,31,31,3,3,3,3,3,3,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{0,0,0,0,0,0,33,1,16,16,16,3,16,16,0,0,0,0,0,3,16,1,16,16,3,16,16,3,16,16,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}};
	end
	
	// Samus Combinational Logic:
	always_comb begin
	   // Determine the width and height of the
		// Defaults:
		color = 0;
		draw = 0;
	   case(sprite_num)
		// SAMUS STAND:
		3'b000: begin
			if(vga_x >= sprite_x && vga_x < sprite_x + width1 && vga_y >= sprite_y && vga_y < sprite_y + height1) begin
			// Output the "draw" signal:
			// Make sure that the pointer is inside the sprite:
				if(direction == 1'b0) begin
					if(samus1[vga_y - sprite_y][vga_x - sprite_x] != 0) begin
						draw = 1'b1;
						color = samus1[vga_y - sprite_y][vga_x - sprite_x];
					end
				end
				if(direction == 1'b1) begin
					if(samus1[vga_y - sprite_y][sprite_x + width1 - 1 - vga_x] != 0) begin
						draw = 1'b1;
						color = samus1[vga_y - sprite_y][sprite_x + width1 - 1 - vga_x];
					end
				end
			end
		end
		// SAMUS WALK 1:
		3'b001: begin
			// Output the "draw" signal:
			// Make sure that the pointer is inside the sprite:
			if(vga_x >= sprite_x && vga_x < sprite_x + width2 && vga_y >= sprite_y && vga_y < sprite_y + height2) begin
				// If the color is not pink output draw:
				if(direction == 1'b0) begin
					if(samus2[vga_y - sprite_y][vga_x - sprite_x] != 0) begin
						draw = 1'b1;
						color = samus2[vga_y - sprite_y][vga_x - sprite_x];
					end
				end
				if(direction == 1'b1) begin
					if(samus2[vga_y - sprite_y][sprite_x + width2 - 1 - vga_x] != 0) begin
						draw = 1'b1;
						color = samus2[vga_y - sprite_y][sprite_x + width2 - 1 - vga_x];
					end
				end
			end
		end
		// SAMUS WALK 2:
		3'b010: begin
			// Output the "draw" signal:
			// Make sure that the pointer is inside the sprite:
			if(vga_x >= sprite_x && vga_x < sprite_x + width3 && vga_y >= sprite_y && vga_y < sprite_y + height3) begin
				// If the color is not pink output draw:
				if(direction == 1'b0) begin
					if(samus3[vga_y - sprite_y][vga_x - sprite_x] != 0) begin
						draw = 1'b1;
						color = samus3[vga_y - sprite_y][vga_x - sprite_x];
					end
				end
				if(direction == 1'b1) begin
					if(samus3[vga_y - sprite_y][sprite_x + width3 - 1 - vga_x] != 0) begin
						draw = 1'b1;
						color = samus3[vga_y - sprite_y][sprite_x + width3 - 1 - vga_x];
					end
				end
			end
		end
		// SAMUS WALK 3:
		3'b011: begin
			// Output the "draw" signal:
			// Make sure that the pointer is inside the sprite:
			if(vga_x >= sprite_x && vga_x < sprite_x + width4 && vga_y >= sprite_y && vga_y < sprite_y + height4) begin
				// If the color is not pink output draw:
				if(direction == 1'b0) begin
					if(samus4[vga_y - sprite_y][vga_x - sprite_x] != 0) begin
						draw = 1'b1;
						color = samus4[vga_y - sprite_y][vga_x - sprite_x];
					end
				end
				if(direction == 1'b1) begin
					if(samus4[vga_y - sprite_y][sprite_x + width4 - 1 - vga_x] != 0) begin
						draw = 1'b1;
						color = samus4[vga_y - sprite_y][sprite_x + width4 - 1 - vga_x];
					end
				end
			end
		end
		// SAMUS JUMP UP:
		3'b100: begin
			// Output the "draw" signal:
			// Make sure that the pointer is inside the sprite:
			if(vga_x >= sprite_x && vga_x < sprite_x + width5 && vga_y >= sprite_y && vga_y < sprite_y + height5) begin
				if(direction == 1'b0) begin
					if(samus5[vga_y - sprite_y][vga_x - sprite_x] != 0) begin
						draw = 1'b1;
						color = samus5[vga_y - sprite_y][vga_x - sprite_x];
					end
				end
				if(direction == 1'b1) begin
					if(samus5[vga_y - sprite_y][sprite_x + width5 - 1 - vga_x] != 0) begin
						draw = 1'b1;
						color = samus5[vga_y - sprite_y][sprite_x + width5 - 1 - vga_x];
					end
				end
			end
		end
		// SAMUS JUMP MOVE:
		3'b101: begin
			// Output the "draw" signal:
			// Make sure that the pointer is inside the sprite:
			if(vga_x >= sprite_x && vga_x < sprite_x + width6 && vga_y >= sprite_y && vga_y < sprite_y + height6) begin
				// If the color is not pink output draw:
				if(direction == 1'b0) begin
					if(samus6[vga_y - sprite_y][vga_x - sprite_x] != 0) begin
						draw = 1'b1;
						color = samus6[vga_y - sprite_y][vga_x - sprite_x];
					end
				end
				if(direction == 1'b1) begin
					if(samus6[vga_y - sprite_y][sprite_x + width6 - 1 - vga_x] != 0) begin
						draw = 1'b1;
						color = samus6[vga_y - sprite_y][sprite_x + width6 - 1 - vga_x];
					end
				end
			end
		end
		// SAMUS standing forward:
		3'b110: begin
			// Output the "draw" signal:
			// Make sure that the pointer is inside the sprite:
			if(vga_x >= sprite_x && vga_x < sprite_x + width7 && vga_y >= sprite_y && vga_y < sprite_y + height7) begin
				// If the color is not pink output draw:
				if(direction == 1'b0) begin
					if(samus7[vga_y - sprite_y][vga_x - sprite_x] != 0) begin
						draw = 1'b1;
						color = samus7[vga_y - sprite_y][vga_x - sprite_x];
					end
				end
				if(direction == 1'b1) begin
					if(samus7[vga_y - sprite_y][sprite_x + width7 - 1 - vga_x] != 0) begin
						draw = 1'b1;
						color = samus7[vga_y - sprite_y][sprite_x + width7 - 1 - vga_x];
					end
				end
			end
		end
		default: begin
			if(vga_x >= sprite_x && vga_x < sprite_x + width1 && vga_y >= sprite_y && vga_y < sprite_y + height1) begin
				// If the color is not pink output draw:
				if(direction == 1'b0) begin
					if(samus1[vga_y - sprite_y][vga_x - sprite_x] != 0) begin
						draw = 1'b1;
						color = samus1[vga_y - sprite_y][vga_x - sprite_x];
					end
				end
				if(direction == 1'b1) begin
					if(samus1[vga_y - sprite_y][sprite_x + width1 - 1 - vga_x] != 0) begin
						draw = 1'b1;
						color = samus1[vga_y - sprite_y][sprite_x + width1 - 1 - vga_x];
					end
				end
			end
		end
		endcase
	end
endmodule

///*

//--------------------------------------------------------------------------------------------
// Monster:
//
//		If the vga pixel pointer is within the monster(s), return a proper color:
//		Priority 2
//		
//--------------------------------------------------------------------------------------------
module monster(
	input logic  			enable1, enable2, enable3,
	input logic  [10:0] 	vga_x, vga_y, sprite1_x, sprite1_y, sprite2_x, sprite2_y, sprite3_x, sprite3_y,
	output logic [5:0] 	color,
	output logic 			draw
);
	// Monster Sprites:
	parameter [9:0] height1 = 30;
	parameter [9:0] width1 = 30;
	parameter [9:0] height2 = 30;
	parameter [9:0] width2 = 45;
	parameter [9:0] height3 = 20;
	parameter [9:0] width3 = 30;
	
	int monster1[height1][width1];
	int monster2[height2][width2];
	int monster3[height3][width3];
	
	always_ff begin
		monster1 =   '{'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,28,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,11,20,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,27,28,33,33,33,33,33,33,33,24,27,33,33,33,33,33,33,33,27,28,33,33,33,33,33},
							'{33,33,33,33,33,11,24,33,33,33,33,33,33,33,2,31,33,33,33,33,33,33,28,11,28,33,33,33,33,33},
							'{33,33,33,33,33,30,30,24,28,33,33,33,24,24,18,30,24,28,33,33,33,24,24,30,31,33,33,33,33,33},
							'{33,33,33,33,33,18,30,11,28,33,33,33,11,11,18,30,11,28,33,33,33,11,24,18,31,33,33,33,33,33},
							'{33,33,33,33,33,18,2,18,24,11,33,33,18,18,2,2,18,33,33,24,11,18,18,2,31,33,33,33,33,33},
							'{33,33,33,33,33,18,18,2,30,11,28,33,2,2,2,2,2,31,33,24,11,18,18,18,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,2,2,2,2,2,2,2,2,2,2,2,2,18,18,2,25,33,33,33,33,33,33,33},
							'{33,28,28,33,33,33,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,25,33,33,33,28,28,33,33},
							'{33,24,24,33,33,33,33,2,2,2,2,2,2,2,2,2,2,2,2,2,2,18,25,33,33,33,24,11,33,33},
							'{33,10,30,25,31,24,27,2,2,2,2,2,2,2,18,2,2,2,2,2,2,2,18,25,27,24,30,30,33,33},
							'{33,25,2,2,2,11,24,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,24,11,30,2,33,33},
							'{33,33,33,18,18,30,18,2,2,2,16,33,33,33,33,33,33,33,33,33,33,2,18,2,18,30,31,33,33,33},
							'{33,33,33,25,18,2,2,2,18,18,33,33,33,33,33,33,33,33,33,33,33,18,18,2,18,18,33,33,33,33},
							'{33,33,33,33,33,2,2,2,31,33,33,33,18,18,18,18,18,18,18,33,33,33,33,2,31,33,33,33,33,33},
							'{33,33,33,33,31,2,18,25,33,33,33,28,25,25,2,2,2,18,25,28,28,33,33,25,31,28,33,33,33,33},
							'{33,33,33,18,2,2,25,33,33,33,24,11,33,33,2,2,2,16,33,24,24,33,33,33,27,11,33,33,19,19},
							'{33,33,33,25,30,18,25,33,33,33,24,11,20,27,31,31,31,27,20,11,24,33,33,33,27,24,1,1,31,33},
							'{33,33,33,27,13,2,25,33,33,33,24,11,11,24,33,33,33,24,11,11,11,33,33,33,31,18,30,30,33,33},
							'{33,31,1,33,33,33,16,25,25,25,28,28,28,28,25,31,19,28,28,33,28,25,25,18,31,33,33,33,33,33},
							'{33,1,30,33,33,33,33,2,2,2,33,33,33,33,2,18,27,33,33,33,33,2,2,2,31,33,33,33,33,33},
							'{33,1,19,33,33,33,33,13,28,33,33,33,33,33,33,31,19,33,33,33,33,33,33,27,1,33,33,33,33,33},
							'{33,1,27,33,33,33,33,19,31,33,33,33,33,33,33,33,19,33,33,33,33,33,33,19,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,19,1,33,24,11,33,33,33,33,33,33,33,24,24,33,33,33,1,27,13,19,33,33},
							'{33,33,33,33,33,33,33,1,28,1,27,20,28,28,33,33,33,28,28,24,20,33,33,33,33,1,1,27,33,33},
							'{33,33,33,33,33,33,33,33,1,27,33,33,11,24,33,33,33,24,11,33,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,28,33,33,28,28,33,33,33,33,28,33,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33}};
							
	   monster2 =   '{'{33,33,33,33,33,33,33,33,33,33,28,27,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,27,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,27,11,28,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,28,11,28,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,24,24,11,24,24,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,24,24,11,24,24,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,28,11,11,11,11,11,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,11,11,11,11,11,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,28,11,24,26,24,11,11,24,33,33,33,33,33,33,33,33,33,33,33,33,33,33,24,11,11,24,26,24,11,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,28,11,24,26,24,11,11,24,33,33,33,33,33,33,33,33,33,33,33,33,33,33,11,11,24,24,26,24,11,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,28,11,24,26,26,26,11,24,33,33,33,33,33,33,33,33,33,33,33,33,33,33,11,24,26,26,26,24,11,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,24,24,24,24,24,24,27,33,33,33,33,33,33,33,33,33,33,33,33,33,5,20,24,24,24,24,24,20,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,27,11,11,11,33,33,23,37,33,33,33,33,33,33,33,33,33,33,37,23,33,28,11,11,11,28,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,37,28,28,28,28,37,37,23,37,33,33,33,33,33,33,33,33,33,33,37,23,37,23,28,28,28,5,37,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,23,37,33,33,33,23,23,23,37,33,33,33,33,33,33,33,33,33,33,37,23,23,37,33,33,33,37,23,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,23,37,37,37,23,23,37,33,33,33,33,33,33,33,33,33,33,33,33,33,33,23,23,37,37,37,23,23,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,23,23,23,23,23,23,37,33,33,33,33,33,33,33,33,33,33,33,33,33,33,23,23,23,23,23,23,23,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,33,37,23,23,23,23,23,23,16,33,33,33,33,33,33,37,37,23,23,23,23,23,37,33,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,16,33,37,37,37,37,37,37,37,16,33,33,33,33,33,33,37,37,37,37,37,37,37,16,16,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,23,23,23,23,23,33,33,33,33,33,33,33,37,23,23,23,23,23,23,16,33,33,33,33,33,33,37,37,23,23,23,23,33,33,33,33,33,33},
							'{33,33,33,33,37,37,37,23,23,23,37,37,33,33,33,33,33,33,37,10,26,23,23,23,23,23,37,37,33,33,33,33,33,33,37,37,23,23,23,37,16,23,33,33,33},
							'{33,33,33,37,37,23,23,23,23,23,16,33,33,33,33,33,33,16,37,24,11,37,23,23,23,23,23,23,33,33,33,33,33,33,33,37,23,23,23,23,23,23,16,33,33},
							'{33,33,37,26,24,23,23,23,23,23,23,37,37,37,33,33,37,37,23,23,23,23,23,23,23,23,23,23,37,37,33,33,37,37,37,23,35,23,23,23,23,24,23,37,33},
							'{33,16,23,26,11,23,23,23,23,23,23,23,23,23,33,33,23,23,23,23,23,23,23,23,23,23,23,23,23,23,33,33,23,23,23,23,23,23,23,23,23,11,26,23,33},
							'{33,23,23,24,11,23,23,23,23,23,23,23,23,23,23,37,33,33,33,37,23,23,23,23,23,23,37,33,33,33,23,23,23,23,23,23,23,23,23,23,23,11,26,23,33},
							'{33,16,23,26,24,23,23,37,37,37,23,23,37,37,23,37,33,33,33,37,37,23,23,23,23,37,16,33,33,33,23,23,37,23,23,37,37,37,37,23,23,24,26,23,33},
							'{33,23,23,23,23,23,23,33,33,33,37,23,16,33,23,23,11,11,11,28,33,37,23,23,37,33,27,11,11,11,37,37,33,16,23,16,33,33,33,23,23,23,23,23,33},
							'{33,33,26,23,23,37,16,33,33,16,37,23,33,33,37,37,11,11,11,24,28,37,37,37,16,27,24,11,11,11,23,16,33,37,23,37,16,33,33,37,37,23,23,26,33},
							'{33,28,11,23,23,33,33,33,33,23,23,23,33,33,33,33,11,11,11,11,11,33,33,33,28,11,11,11,11,11,33,33,33,16,23,23,23,33,33,33,16,23,26,24,28},
							'{33,28,11,24,24,33,33,33,33,26,37,16,33,33,33,33,28,24,11,20,28,37,37,37,5,28,24,11,20,28,33,33,33,33,16,27,26,33,33,33,33,24,24,11,28},
							'{33,28,11,11,11,33,33,33,28,11,27,33,33,33,33,33,33,28,11,28,33,37,23,23,37,33,20,11,28,33,33,33,33,33,33,24,11,33,33,33,28,11,11,11,33},
							'{33,33,33,24,11,33,33,33,33,33,33,33,33,33,33,33,33,33,33,37,37,23,23,23,23,37,23,33,33,33,33,33,33,33,33,33,33,33,33,33,28,11,20,33,33},
							'{33,33,33,20,24,33,33,33,33,33,33,33,33,33,33,33,33,33,33,37,37,23,23,23,23,35,23,33,33,33,33,33,33,33,33,33,33,33,33,33,28,24,27,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33}};

		monster3 = 	 '{'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,3,3,21,3,21,3,21,3,21,33,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,3,21,21,21,21,21,21,21,21,33,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,16,21,21,21,21,21,21,21,21,21,21,21,21,21,21,22,31,33,30,22,33,33},
							'{33,33,33,33,33,33,16,33,16,3,21,21,21,21,21,21,21,21,21,21,21,21,2,22,30,31,25,30,33,33},
							'{33,33,33,33,33,21,21,0,32,33,3,21,21,21,21,21,21,18,22,21,21,22,22,22,22,22,33,33,33,33},
							'{33,33,33,16,16,21,21,21,15,10,16,16,21,21,21,21,2,2,18,16,16,2,7,22,22,18,33,33,31,31},
							'{33,33,33,3,21,21,21,21,21,0,33,33,21,21,21,21,22,18,21,33,33,0,0,22,2,21,33,33,22,22},
							'{33,16,3,16,33,33,33,33,3,21,33,33,21,21,21,21,21,16,33,18,30,21,2,22,22,2,22,22,21,25},
							'{33,16,21,33,33,33,33,33,16,21,33,33,21,21,21,21,21,16,33,22,22,21,18,22,22,22,22,22,21,3},
							'{33,33,33,15,0,0,0,0,32,33,33,33,21,21,21,3,33,25,22,22,22,22,22,22,22,22,21,21,33,33},
							'{33,33,33,0,0,0,0,0,10,33,33,33,3,3,21,3,33,18,22,22,22,22,22,22,22,22,18,21,33,33},
							'{33,10,0,22,22,22,22,0,0,0,21,21,33,16,21,21,21,21,21,22,22,22,22,22,10,33,22,22,22,22},
							'{33,10,0,30,10,10,30,10,15,21,21,21,32,16,16,3,21,21,21,18,2,10,22,22,30,31,10,25,10,31},
							'{33,10,0,33,33,33,33,33,16,21,21,21,0,15,33,16,21,21,21,21,21,33,31,22,22,22,33,33,33,33},
							'{33,33,32,33,33,33,33,33,33,16,16,33,16,33,33,33,16,16,16,33,16,33,33,31,31,31,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33}};
	end
	
	// Monster Combinational Logic:
	always_comb begin
	   // Defaults:
		draw = 0;
		color = 0;
		// Make sure that the pointer is inside the MONSTER 1:
		if(vga_x >= sprite1_x && vga_x < sprite1_x + width1 && vga_y >= sprite1_y && vga_y < sprite1_y + height1 && enable1) begin
		   // If the color is not pink output draw:
			if(monster1[vga_y - sprite1_y][vga_x - sprite1_x] != 33) begin
				draw = 1'b1;
				color = monster1[vga_y - sprite1_y][vga_x - sprite1_x];
			end
		end
		// MONSTER 2
		if(vga_x >= sprite2_x && vga_x < sprite2_x + width2 && vga_y >= sprite2_y && vga_y < sprite2_y + height2 && enable2) begin
		   // If the color is not pink output draw:
			if(monster1[vga_y - sprite2_y][vga_x - sprite2_x] != 33) begin
				draw = 1'b1;
				color = monster2[vga_y - sprite2_y][vga_x - sprite2_x];
			end
		end
		// MONSTER 3
		if(vga_x >= sprite3_x && vga_x < sprite3_x + width3 && vga_y >= sprite3_y && vga_y < sprite3_y + height3 && enable3) begin
		   // If the color is not pink output draw:
			if(monster3[vga_y - sprite3_y][vga_x - sprite3_x] != 33) begin
				draw = 1'b1;
				color = monster3[vga_y - sprite3_y][vga_x - sprite3_x];
			end
		end
	end
endmodule
//*/
/*
//--------------------------------------------------------------------------------------------
// PowerUp:
//
//		If the vga pixel pointer is within the powerUp, return a proper color:
//		Priority 3
//		
//--------------------------------------------------------------------------------------------
module power_up(
	input logic  			enable1, enable2, enable3,
	input logic  [10:0] 	vga_x, vga_y, sprite1_x, sprite1_y, sprite2_x, sprite2_y, sprite3_x, sprite3_y,
	input logic  [1:0] 	sprite_num,
	output logic [5:0] 	color,
	output logic 			draw
);
// Mux the certain power up:
// powerUp Sprites:
	parameter [9:0] height = 70;
	parameter [9:0] width = 45;
	
	int EN[height][width];
	
	always_ff begin
		EN = '{'{33,24,24,24,24,24,24,24,24,24,24,24,24,34,33,29,24,24,29,33,33,33,33,33,29,24,24,34,33},33,
				 '{33,24,24,24,29,29,29,29,29,29,29,29,29,28,33,29,24,24,29,28,33,33,33,33,24,24,24,28,33,33},
				 '{33,24,29,24,29,34,9,29,9,9,9,29,9,5,33,29,24,24,24,24,28,33,33,33,29,24,24,29,33,33},
				 '{33,24,24,24,29,33,33,33,33,33,33,33,33,33,33,29,24,24,24,24,29,28,33,33,29,24,24,28,33,33},
				 '{33,24,24,24,28,33,33,33,33,33,33,33,33,33,33,29,24,24,24,24,24,24,28,33,24,24,24,29,33,33},
				 '{33,24,24,24,29,24,29,24,29,24,29,28,33,33,33,29,24,24,24,24,24,24,29,24,29,24,24,28,33,33},
				 '{33,24,29,24,24,24,29,24,24,29,24,29,33,33,33,29,24,24,29,24,29,24,24,24,24,24,24,34,33,33},
				 '{33,24,24,24,29,9,34,9,9,29,9,5,33,33,33,29,24,24,29,29,29,24,24,24,24,24,24,28,33,33},
				 '{33,24,24,24,29,34,5,37,5,5,34,33,33,33,33,29,24,24,29,34,34,29,24,24,24,24,24,29,33,33},
				 '{33,24,24,24,28,33,33,33,33,33,33,33,33,33,33,29,24,24,29,33,33,9,29,24,24,29,24,28,33,33},
				 '{33,24,29,24,29,28,28,34,28,28,28,34,28,33,33,29,24,24,29,33,33,5,34,29,24,24,24,29,33,33},
				 '{33,24,24,24,24,24,24,24,24,24,24,24,24,34,33,29,24,24,29,33,33,33,5,9,24,24,24,28,33,33},
				 '{33,34,34,29,34,34,29,34,34,34,29,34,29,33,33,34,29,34,34,33,33,33,33,33,34,34,29,34,33,33},
				 '{33,9,23,9,23,9,37,23,9,23,9,37,9,5,33,5,37,9,9,33,33,33,33,33,9,37,9,5,33,33},
				 '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33}};
	end
	
	// Monster Combinational Logic:
	always_comb begin
	   // Defaults:
		draw = 0;
		color = 0;
		// Make sure that the pointer is inside the powerUp 1:
		if(vga_x >= sprite1_x && vga_x < sprite1_x + width && vga_y >= sprite1_y && vga_y < sprite1_y + height && enable1) begin
		   // If the color is not pink output draw:
			//if( != 63)
			draw = 1'b1;
			color = 6'b0;
		end
		// powerUp 2
		if(vga_x >= sprite2_x && vga_x < sprite2_x + width && vga_y >= sprite2_y && vga_y < sprite2_y + height && enable2) begin
		   // If the color is not pink output draw:
			//if( != 63)
			draw = 1'b1;
			color = 6'b0;
		end
		// powerUp 3
		if(vga_x >= sprite3_x && vga_x < sprite3_x + width && vga_y >= sprite3_y && vga_y < sprite3_y + height && enable3) begin
		   // If the color is not pink output draw:
			//if( != 63)
			draw = 1'b1;
			color = 6'b0;
		end
	end
endmodule
*/
///*
//--------------------------------------------------------------------------------------------
// Bullet:
//
//		If the vga pixel pointer is within the bullet(s), return a proper color:
//		Priority 4
//		
//--------------------------------------------------------------------------------------------
module bullet(
	input logic  			enable1, enable2, enable3,
	input logic  [10:0] 	vga_x, vga_y, sprite1_x, sprite1_y, sprite2_x, sprite2_y, sprite3_x, sprite3_y,
	input logic empowered,
	output logic [5:0] 	color,
	output logic 			draw
);
// Mux the bullet instances:
// powerUp Sprites:
	parameter [9:0] height = 10;
	parameter [9:0] width = 10;
	
	int BulletN [height][width];
	int BulletE [height][width];
	
	always_ff begin
	    BulletN = '{'{00,00,00,00,18,18,00,00,00,00},
		             '{00,00,18,18,20,20,18,18,00,00},
						 '{00,18,20,20,20,20,20,20,18,00},
						 '{00,18,20,20,18,18,20,20,18,00},
						 '{18,20,20,18,18,18,18,20,20,18},
						 '{18,20,20,18,18,18,18,20,20,18},
						 '{00,18,20,20,18,18,20,20,18,00},
						 '{00,18,20,20,20,20,20,20,18,00},
						 '{00,00,18,18,20,20,18,18,00,00},
						 '{00,00,00,00,18,18,00,00,00,00}};
		BulletE = '{'{00,00,00,00,06,06,00,00,00,00},
		            '{00,00,06,06,07,07,06,06,00,00},
						'{00,06,07,07,07,07,07,07,06,00},
						'{00,06,07,07,06,06,07,07,06,00},
						'{06,07,07,06,06,06,06,07,07,06},
						'{06,07,07,06,06,06,06,07,07,06},
						'{00,06,07,07,06,06,07,07,06,00},
						'{00,06,07,07,07,07,07,07,06,00},
						'{00,00,06,06,07,07,06,06,00,00},
						'{00,00,00,00,06,06,00,00,00,00}};
	end
	
	// Monster Combinational Logic:
	always_comb begin
	// Defaults:
	color = 0;
	draw = 0;
		// Make sure that the pointer is inside the normal bullet:
		if(vga_x >= sprite1_x && vga_x < sprite1_x + width && vga_y >= sprite1_y && vga_y < sprite1_y + height && enable1) begin
		   // If the color is not pink output draw:
			if(BulletN[vga_x - sprite1_x][vga_y - sprite1_y] != 0) begin
			    draw = 1'b1;
			    color = BulletN[vga_x - sprite1_x][vga_y - sprite1_y];
				 // Enpowered bullet
				 if(empowered == 1'b1) color = BulletE[vga_x - sprite1_x][vga_y - sprite1_y];
			end
		end
		// bullet 2
		if(vga_x >= sprite2_x && vga_x < sprite2_x + width && vga_y >= sprite2_y && vga_y < sprite2_y + height && enable2) begin
		   // If the color is not pink output draw:
			if(BulletN[vga_x - sprite2_x][vga_y - sprite2_y] != 0) begin
			    draw = 1'b1;
			    color = BulletN[vga_x - sprite2_x][vga_y - sprite2_y];
				 // Empowered bullet
				 if(empowered == 1'b1) color = BulletE[vga_x - sprite2_x][vga_y - sprite2_y];
			end
		end
		// Bullet 3
		if(vga_x >= sprite3_x && vga_x < sprite3_x + width && vga_y >= sprite3_y && vga_y < sprite3_y + height && enable3) begin
		   // If the color is not pink output draw:
			if(BulletN[vga_x - sprite3_x][vga_y - sprite3_y] != 0) begin
			    draw = 1'b1;
			    color = BulletN[vga_x - sprite3_x][vga_y - sprite3_y];
				 // Empowered Bullet:
				 if(empowered == 1'b1) color = BulletE[vga_x - sprite3_x][vga_y - sprite3_y];
			end
		end
	end
endmodule
//*/

//--------------------------------------------------------------------------------------------
// Background:
//
//		If the vga pixel pointer is within the proper background tile, return a proper color:
//		Priority 5
//		
//--------------------------------------------------------------------------------------------
module background(
   input logic  [10:0]	background_start_addr,
	input logic  [9:0] 	vga_x, vga_y,
	output logic [5:0] 	color
);
	// Background Tile sizes:
	parameter [9:0] height = 30;
	parameter [9:0] width = 30;
	parameter [9:0] screenH = 16;
	parameter [9:0] screenW = 22;
	// Combinational math an returns 
	logic [10:0] background_x, background_y; // Normalized background array pointers:
	logic [10:0] tile_x, tile_y; // Normalized tile coordinate pointers:
	
	// Sprites: 8 different backgrounds:
	int BG1 [height][width];
	int BG2 [height][width];
	int BG3 [height][width];
	int BG4 [height][width];
	int BG5 [height][width];
	int BG6 [height][width];
	int BG7 [height][width];
	int BG8 [height][width];
	int dummy [screenH][screenW];
	
	//-------------------------------------------------------------------------------------------------------------
	// Sprite arrays + dummy background array:
	//-------------------------------------------------------------------------------------------------------------
	always_ff begin
		dummy = '{'{1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1},
		          '{1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1},
					 '{1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1},
					 '{1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1},
					 '{1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,7,7,6,0,0,1,1},
					 '{1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,7,7,4,0,0,1,1},
					 '{1,0,0,0,0,0,0,1,2,3,3,0,0,0,0,7,7,5,0,0,1,1},
					 '{1,0,0,0,0,0,0,3,2,2,2,0,0,0,0,0,0,0,0,0,1,1},
					 '{1,0,0,0,0,1,1,1,1,0,3,0,0,0,0,0,0,0,0,0,1,1},
					 '{1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1},
					 '{1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1},
					 '{1,0,0,0,0,0,0,0,0,2,3,0,0,0,0,0,0,0,0,0,1,1},
					 '{1,0,0,0,0,0,0,0,0,2,2,0,0,0,0,0,0,0,0,0,1,1},
					 '{1,0,0,0,0,0,0,0,0,2,2,0,0,0,0,0,0,0,0,0,1,1},
					 '{1,0,0,0,0,0,0,0,0,2,2,2,3,2,1,1,1,1,1,1,1,1},
					 '{1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1}};
		// All Black (08):
		BG1 = '{'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
		        '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33}};
		// BLue_brick1:
		BG2 = '{'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
		        '{33,33,33,33,33,33,33,28,33,28,33,28,33,28,33,28,33,28,33,28,33,28,33,28,33,28,33,33,33,33},
				  '{33,33,33,33,33,28,24,26,24,26,24,26,24,26,24,26,24,26,24,26,24,26,24,26,24,26,26,33,33,33},
				  '{33,33,28,28,28,29,29,29,29,29,29,29,29,29,29,29,29,29,29,29,29,29,29,29,29,29,29,33,33,33},
				  '{33,33,26,24,26,26,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,33,33,33},
				  '{33,33,26,26,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,33,33,33},
				  '{33,33,26,26,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,33,33,33},
				  '{33,33,26,26,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,33,33,33},
				  '{33,33,26,26,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,05,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,28,28,28,28,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,28,24,26,24,26,26,33,33,33},
				  '{33,33,28,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,33,33,33,28,26,26,29,29,34,33,33,33},
              '{33,33,26,24,26,24,26,24,26,24,26,24,26,24,26,24,26,26,33,33,33,28,24,29,34,34,34,33,33,33},
              '{33,33,26,26,29,34,29,34,34,29,34,34,29,34,34,29,34,34,33,33,26,29,34,34,34,34,34,33,33,33},
				  '{33,33,26,26,34,34,34,34,34,34,34,34,34,34,34,34,34,34,33,33,26,26,34,34,34,34,34,33,33,33},
				  '{33,33,26,26,34,34,34,34,34,34,34,34,34,34,34,34,34,34,33,33,24,29,34,34,34,34,34,33,33,33},
				  '{33,33,26,26,34,34,34,34,34,34,34,34,34,34,34,34,5,5,33,33,26,26,34,34,34,34,34,33,33,33},
				  '{33,33,26,26,34,34,34,34,34,34,34,34,34,34,34,34,33,33,33,33,26,26,34,34,34,34,34,33,33,33},
				  '{33,33,28,28,5,33,5,33,5,33,5,33,5,33,5,33,33,33,33,33,28,34,33,5,33,5,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,26,26,26,26,26,26,26,33,33,33,33,33,33,33,33,33,33,33,26,26,26,26,26,26,27,33,33,33},
				  '{33,33,26,24,26,24,26,24,26,33,33,33,33,33,33,33,33,33,33,33,26,24,26,24,26,24,26,33,33,33},
				  '{33,33,26,26,34,34,34,34,34,34,34,34,34,34,34,34,34,34,26,26,34,34,34,34,34,34,34,33,33,33},
				  '{33,33,26,26,34,34,34,34,34,34,34,34,34,34,34,34,34,34,26,26,34,34,34,34,34,34,34,33,33,33},
				  '{33,33,26,26,34,34,34,34,34,34,34,34,34,34,34,34,34,34,24,26,34,34,34,34,34,34,34,33,33,33},
				  '{33,33,28,27,5,5,5,5,5,5,5,5,5,5,5,5,5,5,27,28,5,5,5,5,5,5,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33}};
		
		// Brick grey:
		BG3 =     '{'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,33,33},
						'{33,33,33,33,33,33,10,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,26,33,33},
						'{33,33,33,26,26,26,22,26,30,26,22,30,26,22,30,26,22,30,26,22,30,26,22,30,26,22,30,10,33,33},
						'{33,33,33,7,7,7,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,10,33,33},
						'{33,33,33,7,22,30,30,30,30,30,10,30,30,10,30,30,10,30,30,10,30,30,10,30,30,10,30,10,33,33},
						'{33,33,33,7,7,10,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,10,33,33},
						'{33,33,33,7,7,10,30,30,30,10,30,10,30,30,10,30,30,10,30,30,10,30,30,10,30,30,30,10,33,33},
						'{33,33,33,10,10,32,32,31,32,32,31,10,31,32,31,32,31,32,31,32,31,32,31,32,31,32,31,31,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,32,30,30,30,30,10,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,10,7,7,7,7,26,33,33},
						'{33,33,33,26,22,26,7,26,22,26,7,26,22,26,7,26,22,26,22,33,33,33,10,7,26,30,30,10,33,33},
						'{33,33,33,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,26,33,33,33,10,7,30,30,30,10,33,33},
						'{33,33,33,7,7,10,30,30,10,30,30,10,30,30,10,30,30,30,10,33,31,7,26,30,30,30,30,10,33,33},
						'{33,33,33,7,22,30,30,30,30,30,30,30,30,30,30,30,10,30,10,33,32,7,22,30,30,30,30,10,33,33},
						'{33,33,33,7,7,10,30,30,30,10,30,10,30,10,30,30,30,30,10,33,32,7,26,30,30,10,30,10,33,33},
						'{33,33,33,7,26,30,30,30,30,30,30,30,30,30,10,30,10,31,33,33,32,7,22,30,30,30,30,10,33,33},
						'{33,33,33,7,7,10,30,10,30,10,30,30,10,30,30,30,30,33,33,33,32,7,26,30,30,30,30,10,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,7,7,7,7,7,7,7,33,33,33,33,33,33,33,33,33,33,31,7,7,7,7,7,7,26,33,33},
						'{33,33,33,7,7,7,7,7,7,26,33,33,33,33,33,33,33,33,33,33,10,7,7,7,7,7,22,26,33,33},
						'{33,33,33,7,7,10,10,30,30,30,30,30,30,30,30,30,30,30,30,7,7,10,10,10,10,10,30,10,33,33},
						'{33,33,33,7,22,10,30,30,30,30,30,30,30,30,30,30,30,30,30,7,26,30,30,30,30,30,30,10,33,33},
						'{33,33,33,7,7,10,30,30,30,30,30,30,10,30,10,30,10,30,30,7,22,30,30,30,30,10,30,10,33,33},
						'{33,33,33,32,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,32,32,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33}};
		// Brick green:
		BG4 =     '{'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,31,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,33,33,33},
						'{33,33,33,33,33,31,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,25,33,33,33},
						'{33,33,18,18,18,13,20,19,19,20,19,19,19,19,19,19,19,19,19,20,19,19,19,19,20,19,20,33,33,33},
						'{33,33,18,18,25,27,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,33,33,33},
						'{33,33,18,18,19,20,20,19,20,19,20,19,20,19,20,19,20,20,19,20,19,20,20,19,20,20,20,33,33,33},
						'{33,33,18,18,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,19,20,20,19,20,20,33,33,33},
						'{33,33,18,18,19,20,20,19,20,19,20,19,20,19,20,20,20,19,20,19,20,20,20,19,20,20,20,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,31,18,18,18,18,18,33,33,33},
						'{33,33,33,16,33,31,33,16,33,31,33,16,33,31,33,16,33,31,33,33,33,31,18,18,13,18,25,33,33,33},
						'{33,33,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,33,33,33,31,18,19,20,20,20,33,33,33},
						'{33,33,18,18,13,27,25,13,27,25,13,27,25,27,13,25,27,25,33,33,31,25,25,19,20,19,20,33,33,33},
						'{33,33,18,18,20,20,20,20,20,20,20,20,19,20,20,20,19,20,33,33,18,13,20,20,20,20,20,33,33,33},
						'{33,33,18,18,19,20,19,20,19,20,19,20,20,20,19,20,20,20,33,33,18,25,19,20,19,20,20,33,33,33},
						'{33,33,18,18,19,20,20,20,20,20,20,20,20,20,20,19,20,20,33,33,18,13,20,20,20,20,20,33,33,33},
						'{33,33,18,18,19,20,19,20,19,20,20,20,19,20,20,20,33,33,33,33,18,25,19,20,19,20,20,33,33,33},
						'{33,33,25,25,20,28,20,27,20,27,20,27,20,27,20,20,33,33,33,33,18,31,20,28,20,28,28,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,31,31,31,31,31,31,31,33,33,33,33,33,33,33,33,33,33,33,31,31,31,31,31,31,31,33,33,33},
						'{33,33,18,18,18,18,18,18,18,33,33,33,33,33,33,33,33,33,33,33,18,18,18,18,18,18,18,33,33,33},
						'{33,33,18,18,19,27,19,27,19,28,28,28,28,28,28,28,28,28,25,25,27,19,27,19,27,19,27,33,33,33},
						'{33,33,18,18,19,20,20,20,20,19,20,19,19,20,19,19,20,19,18,18,20,20,20,20,20,20,20,33,33,33},
						'{33,33,18,18,20,20,19,20,20,20,20,20,20,20,20,20,20,20,18,18,19,20,20,19,20,20,20,33,33,33},
						'{33,33,18,25,20,20,20,20,20,20,20,20,20,20,20,20,20,20,18,25,20,20,20,20,20,20,28,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33}};
		// Blue door bot mid 1:
		BG5 =     '{'{3,34,29,29,34,29,34,29,34,29,34,29,34,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{2,29,29,29,29,29,29,29,29,29,29,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{25,29,34,29,29,34,29,29,34,29,29,29,34,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,34,29,29,29,29,29,29,29,29,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,29,34,29,34,29,34,29,29,29,29,29,29,34,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,34,29,29,29,29,29,29,34,29,34,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,29,34,29,29,29,34,29,29,29,29,29,34,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,34,29,29,34,29,29,29,29,34,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,29,34,29,29,29,29,34,29,29,29,34,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,34,29,29,29,34,29,29,29,29,29,29,29,34,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,29,34,29,29,29,29,29,34,29,29,34,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,34,29,29,29,34,29,29,29,29,29,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,29,34,29,29,29,29,34,29,34,29,34,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,34,29,29,34,29,29,29,29,29,29,29,29,34,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,29,34,29,29,29,34,29,29,34,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{18,29,29,29,29,29,29,29,29,29,29,34,29,34,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{18,29,34,29,34,29,29,34,29,34,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,34,29,29,29,29,29,29,29,29,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,29,34,29,29,34,29,34,29,29,34,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,29,29,29,29,29,29,29,29,29,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,29,34,29,29,34,29,29,34,29,34,29,34,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,29,29,29,29,29,29,29,29,29,29,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{3,34,29,29,34,29,34,29,34,29,29,34,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,34,29,29,29,29,29,29,29,29,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{3,34,29,34,29,29,34,29,29,34,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,34,29,29,29,29,29,29,29,29,29,34,29,34,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{3,34,29,29,34,29,29,34,29,34,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,34,29,29,29,29,29,29,29,29,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,34,29,29,34,29,34,29,29,34,29,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{21,29,29,29,29,29,29,29,29,29,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}};
		// Blue Door Bot Right:
		BG6 =  '{'{21,29,29,29,29,29,29,29,29,29,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{2,29,34,29,29,34,29,34,29,34,29,29,29,34,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,29,29,29,29,29,29,29,29,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,29,34,29,29,34,29,29,34,29,34,29,34,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,29,29,29,29,29,29,29,29,29,28,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,34,29,34,29,34,29,29,34,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,34,29,29,29,29,29,29,29,29,29,29,5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,29,34,29,29,34,29,29,34,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,34,29,29,29,29,29,29,29,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,34,29,34,29,24,26,29,34,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,34,29,29,29,29,29,26,7,29,29,29,5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,29,29,34,29,26,7,34,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,34,29,29,29,29,24,26,26,29,29,34,28,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,34,29,24,7,26,29,29,29,29,5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,29,29,29,29,24,7,29,29,34,29,34,33,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{2,29,29,34,29,34,24,7,26,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,29,29,26,26,7,7,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,34,24,7,7,7,26,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,7,7,7,24,29,29,34,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,29,7,7,7,26,29,29,29,34,28,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,7,7,7,24,34,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,29,7,7,26,26,29,34,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,7,26,34,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,29,24,26,29,29,34,28,5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,34,29,34,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,34,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,28,34,28,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}};
		// Blue Door bottop:
		BG7 =  '{'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{31,28,5,5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{2,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,34,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,34,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,29,29,34,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,29,29,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,7,26,29,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,29,7,26,24,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,7,7,7,24,29,34,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,29,7,7,7,26,29,29,34,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,7,7,7,24,29,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,29,29,24,7,7,7,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,26,7,7,7,26,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,34,29,34,29,24,7,26,34,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,29,29,29,34,24,7,26,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{2,29,34,29,29,29,24,7,29,29,29,34,29,5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{25,34,29,29,34,29,26,26,24,24,34,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,29,29,29,29,26,7,29,29,29,5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,34,29,29,34,29,29,26,7,29,34,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,29,29,29,29,26,7,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,34,29,29,34,29,29,29,34,29,29,34,28,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,29,29,34,29,29,29,29,29,34,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,34,29,34,29,29,29,34,29,34,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,29,29,29,29,29,29,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,34,29,29,34,29,34,29,29,34,29,34,28,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,29,29,29,29,29,29,29,29,29,34,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,34,29,29,34,29,29,34,29,29,34,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,29,29,29,29,29,29,29,29,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{3,34,29,29,34,29,34,29,34,29,34,29,34,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}};
		// Blue Door left:
		BG8 =  '{'{33,21,21,21,25,21,21,25,21,21,25,21,21,21,21,21,21,21,21,25,21,21,25,21,21,21,25,21,21,29},
					'{16,18,2,2,2,2,2,2,2,2,2,2,2,18,2,18,2,18,2,2,2,2,2,2,2,2,2,2,2,29},
					'{33,2,10,29,24,29,24,29,29,24,29,24,29,16,16,2,30,29,24,29,29,24,29,24,29,29,24,32,16,29},
					'{16,2,24,29,29,29,29,29,29,29,29,29,24,16,16,2,30,29,29,29,29,29,29,29,29,24,29,33,16,29},
					'{33,2,10,29,33,16,16,16,16,16,16,28,29,16,16,18,30,29,28,16,16,16,16,16,16,28,29,28,16,34},
					'{16,2,24,29,16,16,32,33,32,16,16,26,29,16,16,2,30,29,28,16,16,28,32,16,16,10,24,33,16,34},
					'{33,2,24,29,33,16,29,29,24,26,2,24,29,16,16,2,30,29,28,16,29,29,29,24,2,10,29,28,16,29},
					'{16,2,10,29,16,16,29,24,29,24,2,24,29,16,16,2,10,29,28,16,29,24,29,24,18,10,29,31,16,34},
					'{33,2,24,29,33,16,29,29,24,26,2,24,29,16,16,2,30,29,28,16,28,29,29,24,18,10,24,28,16,29},
					'{16,2,24,29,16,16,30,30,30,18,2,26,29,16,16,2,30,29,28,16,25,30,30,18,2,26,29,28,16,34},
					'{33,2,10,29,28,16,2,18,2,2,2,24,29,16,16,2,10,29,28,16,2,2,2,2,2,10,29,28,16,29},
					'{16,2,24,29,29,24,29,29,29,24,29,29,24,16,16,2,30,29,24,29,29,29,29,24,29,24,29,28,16,34},
					'{33,18,10,29,29,28,29,29,29,28,29,29,29,16,16,18,25,29,29,29,29,27,29,29,29,34,29,16,16,29},
					'{33,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,34},
					'{33,21,16,25,16,25,16,25,16,25,16,25,3,25,21,16,25,3,25,16,25,16,25,3,25,16,25,21,16,29},
					'{33,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,18,2,2,29},
					'{16,2,10,26,26,24,26,24,26,24,26,24,26,25,16,2,18,24,26,24,26,24,26,24,26,24,24,10,16,29},
					'{33,2,10,29,24,29,29,29,24,29,29,29,24,16,3,2,30,29,29,24,29,29,29,24,29,29,29,31,16,34},
					'{16,2,24,29,28,16,16,16,16,33,16,29,29,16,16,18,30,29,28,16,33,16,16,16,33,28,29,28,16,34},
					'{33,2,24,29,16,16,16,16,16,16,16,28,29,16,16,2,30,29,28,16,16,16,16,16,3,32,29,31,16,29},
					'{16,2,10,29,33,16,29,29,24,26,2,24,29,16,16,2,10,29,28,16,29,29,29,24,18,10,24,28,16,34},
					'{33,2,24,29,16,16,24,29,29,24,2,26,29,16,16,2,30,29,28,16,29,24,29,24,2,26,29,28,16,29},
					'{16,2,24,29,28,16,29,24,29,24,2,24,29,16,16,2,30,29,28,16,28,29,24,29,2,10,29,28,16,34},
					'{33,2,10,29,16,16,10,26,10,30,18,24,29,16,16,2,10,29,28,16,10,10,26,10,2,10,24,28,16,29},
					'{16,2,24,29,33,16,2,2,2,2,2,26,29,16,16,2,30,29,28,16,21,2,2,2,2,10,29,28,16,34},
					'{33,2,24,29,29,29,26,24,26,26,24,29,24,16,16,18,30,29,29,29,26,24,26,24,29,24,29,28,16,29},
					'{16,2,10,29,24,29,29,29,24,29,29,24,29,16,16,2,10,24,29,24,29,29,29,24,29,29,24,33,16,34},
					'{33,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,29},
					'{33,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,34},
					'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33}};
	end
	
	
	always_comb begin
		// Determines the upper left corner of the tile sprite:
		// Defaults:
		background_x = 0;
		background_y = 0;
		tile_x = 0;
		tile_y = 0;
		
		if(vga_x >= 0 && vga_x < width) begin
	   	background_x = 0;
			tile_x = 0;
		end
		if(vga_x >= width && vga_x < 2*width) begin
			background_x = width;
			tile_x = 1;
		end
		if(vga_x >= 2*width && vga_x < 3*width) begin
			background_x = 2*width;
			tile_x = 2;
		end
		if(vga_x >= 3*width && vga_x < 4*width) begin
			background_x = 3*width;
			tile_x = 3;
		end
		if(vga_x >= 4*width && vga_x < 5*width) begin 
			background_x = 4*width;
			tile_x = 4;
		end
		if(vga_x >= 5*width && vga_x < 6*width) begin
			background_x = 5*width;
			tile_x = 5;
		end
		if(vga_x >= 6*width && vga_x < 7*width) begin
			background_x = 6*width;
			tile_x = 6;
		end
		if(vga_x >= 7*width && vga_x < 8*width) begin
			background_x = 7*width;
			tile_x = 7;
		end
		if(vga_x >= 8*width && vga_x < 9*width) begin
			background_x = 8*width;
			tile_x = 8;
		end
		if(vga_x >= 9*width && vga_x < 10*width) begin
			background_x = 9*width;
			tile_x = 9;
		end
		if(vga_x >= 10*width && vga_x < 11*width) begin
			background_x = 10*width;
			tile_x = 10;
		end
		if(vga_x >= 11*width && vga_x < 12*width) begin
			background_x = 11*width;
			tile_x = 11;
		end
		if(vga_x >= 12*width && vga_x < 13*width) begin
			background_x = 12*width;
			tile_x = 12;
		end
		if(vga_x >= 13*width && vga_x < 14*width) begin
			background_x = 13*width;
			tile_x = 13;
		end
		if(vga_x >= 14*width && vga_x < 15*width) begin
			background_x = 14*width;
			tile_x = 14;
		end
		if(vga_x >= 15*width && vga_x < 16*width) begin
			background_x = 15*width;
			tile_x = 15;
		end
		if(vga_x >= 16*width && vga_x < 17*width) begin
			background_x = 16*width;
			tile_x = 16;
		end
		if(vga_x >= 17*width && vga_x < 18*width) begin
			background_x = 17*width;
			tile_x = 17;
		end
		if(vga_x >= 18*width && vga_x < 19*width) begin
			background_x = 18*width;
			tile_x = 18;
		end
		if(vga_x >= 19*width && vga_x < 20*width) begin
			background_x = 19*width;
			tile_x = 19;
		end
		if(vga_x >= 20*width && vga_x < 21*width) begin
			background_x = 20*width;
			tile_x = 20;
		end
		if(vga_x >= 21*width && vga_x < 22*width) begin
			background_x = 21*width;
			tile_x = 21;
		end
		
		
		if(vga_y >= 0 && vga_y < height) begin
			background_y = 0;
			tile_y = 0;
		end
		if(vga_y >= height && vga_y < 2*height) begin
			background_y = height;
			tile_y = 1;
		end
		if(vga_y >= 2*height && vga_y < 3*height) begin
			background_y = 2*height;
			tile_y = 2;
		end
		if(vga_y >= 3*height && vga_y < 4*height) begin
			background_y = 3*height;
			tile_y = 3;
		end
		if(vga_y >= 4*height && vga_y < 5*height) begin
			background_y = 4*height;
			tile_y = 4;
		end
		if(vga_y >= 5*height && vga_y	< 6*height) begin
			background_y = 5*height;
			tile_y = 5;
		end
		if(vga_y >= 6*height && vga_y < 7*height) begin
			background_y = 6*height;
			tile_y = 6;
		end
		if(vga_y >= 7*height && vga_y < 8*height) begin
			background_y = 7*height;
			tile_y = 7;
		end
		if(vga_y >= 8*height && vga_y < 9*height) begin
			background_y = 8*height;
			tile_y = 8;
		end
		if(vga_y >= 9*height && vga_y < 10*height) begin
			background_y = 9*height;
			tile_y = 9;
		end
		if(vga_y >= 10*height && vga_y < 11*height) begin
			background_y = 10*height;
			tile_y = 10;
		end
		if(vga_y >= 11*height && vga_y < 12*height) begin
			background_y = 11*height;
			tile_y = 11;
		end
		if(vga_y >= 12*height && vga_y < 13*height) begin
			background_y = 12*height;
			tile_y = 12;
		end
		if(vga_y >= 13*height && vga_y < 14*height) begin
			background_y = 13*height;
			tile_y = 13;
		end
		if(vga_y >= 14*height && vga_y < 15*height) begin
			background_y = 14*height;
			tile_y = 14;
		end
		if(vga_y >= 15*height && vga_y < 16*height) begin
			background_y = 15*height;
			tile_y = 15;
		end
	end
	
	// Select the correct background tile from the background tile array:
	always_comb begin
		 // Default == Black
		 color = 33;
		 case(dummy[tile_y][tile_x])
			 0: begin
				color = BG1[vga_y - background_y][vga_x - background_x];
			 end
			 1: begin
				color = BG2[vga_y - background_y][vga_x - background_x];
			 end
			 2: begin
				color = BG3[vga_y - background_y][vga_x - background_x];
			 end
			 3: begin
				color = BG4[vga_y - background_y][vga_x - background_x];
			 end
			 4: begin
				color = BG5[vga_y - background_y][vga_x - background_x];
			 end
			 5: begin
				color = BG6[vga_y - background_y][vga_x - background_x];
			 end
			 6: begin
				color = BG7[vga_y - background_y][vga_x - background_x];
			 end
			 7: begin
				color = BG8[vga_y - background_y][vga_x - background_x];
			 end
			 default: begin
				color = 8;
			 end
		 endcase
		 if(color == 0) color = 33;
	end
endmodule

//
// Controls the title 
module gui(
   input logic titleEn,
	input logic [1:0] health,
	input logic [9:0] vga_x, vga_y,
	output logic [5:0] color,
	output logic draw
);

	// Health Sprites:
	parameter height1 = 15;
	parameter width1 = 30;
	
	parameter height2 = 8;
	parameter width2 = 8;
	
	parameter en_x = 20;
	parameter en_y = 20;
	parameter health1_x = 55;
	parameter health2_x = 65;
	parameter health3_x = 75;
	parameter health_y = 23;
	
	int EN[height1][width1];
	int EN_indicator[height2][width2];
	
	always_ff begin
		EN = '{'{33,24,24,24,24,24,24,24,24,24,24,24,24,34,33,29,24,24,29,33,33,33,33,33,29,24,24,34,33,33},
				 '{33,24,24,24,29,29,29,29,29,29,29,29,29,28,33,29,24,24,29,28,33,33,33,33,24,24,24,28,33,33},
				 '{33,24,29,24,29,34,9,29,9,9,9,29,9,5,33,29,24,24,24,24,28,33,33,33,29,24,24,29,33,33},
				 '{33,24,24,24,29,33,33,33,33,33,33,33,33,33,33,29,24,24,24,24,29,28,33,33,29,24,24,28,33,33},
				 '{33,24,24,24,28,33,33,33,33,33,33,33,33,33,33,29,24,24,24,24,24,24,28,33,24,24,24,29,33,33},
				 '{33,24,24,24,29,24,29,24,29,24,29,28,33,33,33,29,24,24,24,24,24,24,29,24,29,24,24,28,33,33},
				 '{33,24,29,24,24,24,29,24,24,29,24,29,33,33,33,29,24,24,29,24,29,24,24,24,24,24,24,34,33,33},
				 '{33,24,24,24,29,9,34,9,9,29,9,5,33,33,33,29,24,24,29,29,29,24,24,24,24,24,24,28,33,33},
				 '{33,24,24,24,29,34,5,37,5,5,34,33,33,33,33,29,24,24,29,34,34,29,24,24,24,24,24,29,33,33},
				 '{33,24,24,24,28,33,33,33,33,33,33,33,33,33,33,29,24,24,29,33,33,9,29,24,24,29,24,28,33,33},
				 '{33,24,29,24,29,28,28,34,28,28,28,34,28,33,33,29,24,24,29,33,33,5,34,29,24,24,24,29,33,33},
				 '{33,24,24,24,24,24,24,24,24,24,24,24,24,34,33,29,24,24,29,33,33,33,5,9,24,24,24,28,33,33},
				 '{33,34,34,29,34,34,29,34,34,34,29,34,29,33,33,34,29,34,34,33,33,33,33,33,34,34,29,34,33,33},
				 '{33,9,23,9,23,9,37,23,9,23,9,37,9,5,33,5,37,9,9,33,33,33,33,33,9,37,9,5,33,33},
				 '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33}};
		
		EN_indicator =  '{'{33,33,33,33,33,33,33,33},
								'{33,33,25,18,18,25,33,33},
								'{33,33,25,2,18,18,33,33},
								'{33,33,25,2,2,25,33,33},
								'{33,33,25,21,21,25,33,33},
								'{33,33,16,3,3,3,33,33},
								'{33,33,33,16,16,33,33,33},
								'{33,33,33,33,33,33,33,33}};		 
	end
	
	always_comb begin
	   // Defaults:
	   color = 0;
	   draw = 0;
	   
		// Always show the energy:
		if(vga_x >= en_x && vga_x < en_x + width1 && vga_y >= en_y && vga_y < en_y + height1) begin
		   // If the color is not pink output draw:
			if(EN[vga_y - en_x][vga_x - en_x] != 33) begin
			    draw = 1'b1;
			    color = EN[vga_y - en_y][vga_x - en_x];
			end
		end
		// *
		if(vga_x >= health1_x && vga_x < health1_x + width2 && vga_y >= health_y && vga_y < health_y + height2 && (health >= 2'b01)) begin
		   // If the color is not pink output draw:
			if(EN_indicator[vga_y - health_y][vga_x - health1_x] != 33) begin
			    draw = 1'b1;
			    color = EN_indicator[vga_y - health_y][vga_x - health1_x];
			end
		end
		// **
		if(vga_x >= health2_x && vga_x < health2_x + width2 && vga_y >= health_y && vga_y < health_y + height2 && (health >= 2'b10)) begin
		   // If the color is not pink output draw:
			if(EN_indicator[vga_y - health_y][vga_x - health2_x] != 0) begin
			    draw = 1'b1;
			    color = EN_indicator[vga_y - health_y][vga_x - health2_x];
			end
		end
		// ***
		if(vga_x >= health3_x && vga_x < health3_x + width2 && vga_y >= health_y && vga_y < health_y + height2 && (health >= 2'b11)) begin
		   // If the color is not pink output draw:
			if(EN_indicator[vga_y - health_y][vga_x - health3_x] != 33) begin
			    draw = 1'b1;
			    color = EN_indicator[vga_y - health_y][vga_x - health3_x];
			end
		end
	end
endmodule

//--------------------------------------------------------------------------------------------
// Explosions:
//
//		If a monster is destroyed, display the explosions:
//		
//--------------------------------------------------------------------------------------------
module explosion(
	input logic enable1, enable2, enable3, vsync, 
	input logic [9:0] vga_x, vga_y, exp1_x, exp1_y, exp2_x, exp2_y, exp3_x, exp3_y,
	output logic [5:0] color,
	output logic draw
);
	//Sprites:
	parameter height1 = 60;
	parameter width1 = 60;
	
	parameter height2 = 60;
	parameter width2 = 60;
	
	int explosion1[height1][width1];
	int explosion2[height2][width2];
	
	logic vsync_slow[3:0];
	logic [1:0] counter1, counter2, counter3;
	logic released1, released2, released3;
	
	 always_ff @ (posedge vsync)
    begin 
            vsync_slow[0] <= ~ (vsync_slow[0]);
    end
	 always_ff @ (posedge vsync_slow[0])
    begin 
            vsync_slow[1] <= ~ (vsync_slow[1]);
    end
	 always_ff @ (posedge vsync_slow[1])
    begin 
            vsync_slow[2] <= ~ (vsync_slow[2]);
    end
	 always_ff @ (posedge vsync_slow[2])
    begin 
            vsync_slow[3] <= ~ (vsync_slow[3]);
    end

	always_ff begin
		// Small
		explosion1 = '{'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,33,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,33},
							'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,33,33,33,33,8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8,33},
							'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8,33},
							'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8,33},
							'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8,33},
							'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8,33},
							'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8,33},
							'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8,33},
							'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8,33},
							'{8,8,8,8,8,8,8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8,33},
							'{8,8,8,8,8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8,33},
							'{8,8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8,33},
							'{8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8,33},
							'{8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8,8},
							'{8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,21,21,33,33,33,10,0,33,33,33,33,0,32,33,33,33,21,21,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,16,16,33,33,16,10,10,16,16,16,32,10,31,16,33,33,16,16,33,33,33,33,16,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,16,16,33,33,33,33,33,33,16,21,16,33,21,21,21,16,33,16,21,33,33,33,33,33,33,33,16,21,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,10,10,33,33,10,32,33,16,21,15,30,33,16,16,32,30,15,21,33,33,10,32,33,33,30,32,16,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,10,0,33,33,0,30,33,16,21,0,0,33,33,33,33,0,2,21,33,33,0,30,33,32,0,32,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,16,33,15,21,21,0,0,32,33,30,0,21,21,21,15,0,10,33,30,0,21,21,21,31,33,16,21,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,16,16,33,25,21,21,2,0,32,33,30,0,21,21,21,2,0,32,33,30,0,21,2,21,32,33,16,21,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,10,0,19,19,0,30,33,32,0,27,19,0,0,0,26,19,30,0,33,33,0,26,19,27,0,32,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,30,0,19,19,30,10,28,31,0,31,20,30,10,30,10,20,10,0,31,28,10,10,19,30,0,10,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,32,0,0,19,19,33,33,19,25,21,33,33,33,33,33,33,33,16,21,19,19,33,33,19,27,0,0,0,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,32,0,0,30,31,33,33,19,1,16,33,33,28,28,28,28,33,33,16,20,19,33,33,25,18,0,0,0,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,32,0,0,21,21,33,33,19,20,33,33,33,20,19,19,20,33,33,33,20,19,33,33,21,0,0,0,0,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,15,0,0,0,21,21,33,33,19,28,33,33,33,20,19,19,1,33,33,33,20,19,33,33,21,2,0,0,0,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,21,0,0,0,2,21,33,33,19,1,33,33,33,20,19,19,20,33,33,33,20,19,33,33,21,2,0,0,0,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,0,0,0,0,27,19,33,33,19,27,21,33,33,33,33,33,33,33,16,21,19,19,33,33,19,30,0,0,0,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,21,0,0,0,19,19,33,33,20,31,21,31,33,33,33,33,33,33,31,21,1,20,33,33,19,27,0,0,30,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,30,33,32,0,19,19,0,30,33,32,0,27,19,0,0,0,30,19,30,0,28,33,0,26,19,30,0,32,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,10,16,10,10,25,25,0,0,32,10,10,27,30,0,2,0,30,30,10,10,32,32,0,2,25,10,10,32,16,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,21,16,33,16,21,21,21,0,32,33,10,0,21,21,21,0,0,32,33,30,0,21,21,21,16,33,16,21,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,16,32,10,32,16,0,0,32,32,16,0,0,16,16,33,10,0,15,16,10,32,0,0,33,32,30,32,16,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,10,0,33,33,0,30,33,16,21,0,0,33,33,33,32,0,2,21,33,33,0,30,33,32,0,32,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,21,16,33,33,33,33,33,33,16,21,16,33,15,21,21,16,33,16,21,33,33,33,33,33,33,33,16,21,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,21,16,33,33,33,33,33,33,16,21,33,33,21,25,21,16,33,31,21,33,33,33,33,33,33,33,16,21,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,21,21,33,33,33,10,0,33,33,33,28,0,10,33,33,33,21,21,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,16,16,33,33,33,32,30,33,33,33,33,30,28,33,33,33,16,16,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{8,8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{33,8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8},
							'{33,8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8},
							'{33,8,8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8},
							'{33,33,8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8,8,8,8,8,8,8,8,33,33,33,33,33,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8},
							'{33,33,8,8,8,8,8,33,33,33,33,33,33,33,33,33,33,33,33,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,33,33,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8},
							'{33,33,8,8,8,8,8,33,33,33,33,33,33,33,33,33,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8},
							'{33,33,8,8,8,8,8,8,33,33,33,33,33,33,33,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,33,33,33,33,33,33,8,8,8,8,8,8,8},
							'{33,33,8,8,8,8,8,8,33,33,33,33,33,33,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,33,33,33,33,33,33,33,33,8,8,8,8,8,8,8},
							'{8,33,33,8,8,8,8,8,33,33,33,33,33,33,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,33,8,8,8,8,8,8,8},
							'{8,8,33,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8},
							'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8},
							'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8},
							'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8},
							'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8},
							'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8},
							'{8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8}};
		
		// Large
		explosion2 = '{'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,21,16,33,33,33,30,30,33,33,33,32,0,33,33,33,33,21,16,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,21,16,33,33,33,0,30,33,33,33,10,0,33,33,33,33,21,16,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,16,21,33,33,33,33,33,33,33,16,21,33,33,21,21,21,16,33,21,21,33,33,33,33,33,33,33,21,21,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,16,16,32,33,33,33,33,33,33,16,21,32,32,16,25,3,32,33,21,21,33,33,33,33,33,33,33,16,31,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,33,33,0,30,33,33,33,30,0,33,33,0,10,33,16,21,0,0,33,33,33,10,0,21,21,33,33,0,10,33,10,0,33,33,33,28,0,32,33,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,16,16,32,28,33,33,16,10,32,16,10,2,15,10,32,16,0,0,16,16,16,30,0,10,16,10,10,0,15,16,32,10,16,16,33,33,32,32,16,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,21,21,33,33,33,16,21,33,33,21,21,21,2,0,32,33,0,0,21,21,21,0,0,33,33,0,0,21,21,21,16,33,21,21,33,33,33,16,21,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,30,10,33,30,30,19,27,0,10,33,10,30,19,27,0,0,0,30,19,30,30,33,32,0,30,19,10,30,33,33,30,10,33,33,33,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,28,0,32,33,30,0,19,19,0,10,33,30,0,19,19,0,0,0,27,19,26,0,33,33,0,30,19,30,0,33,33,0,30,33,33,33,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,0,10,33,33,33,0,0,33,16,21,0,0,0,0,19,20,33,28,19,25,21,33,33,33,33,33,33,33,21,21,19,20,33,28,19,30,0,0,0,21,16,33,10,0,33,33,33,33,0,10,33,33,33,33},
							'{33,33,33,33,33,33,0,32,33,33,33,30,0,33,33,21,2,0,0,0,19,1,33,28,19,31,21,33,33,33,33,33,33,33,16,25,19,20,33,33,19,26,0,0,0,21,15,33,10,0,33,33,33,33,0,32,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,21,21,33,33,21,0,0,0,0,21,15,33,28,19,28,33,33,33,19,19,19,28,33,33,33,19,20,33,16,21,0,0,0,0,21,16,33,16,21,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,16,33,33,33,16,15,2,32,32,25,2,0,30,30,16,16,33,33,1,33,33,33,33,28,1,1,33,33,33,33,28,28,33,33,16,10,30,0,0,25,10,32,15,0,16,16,33,33,16,33,33,33,33,33},
							'{33,33,33,33,33,33,21,16,33,16,21,0,0,0,30,19,30,0,19,19,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,20,19,0,0,19,27,0,0,0,2,21,33,33,21,16,33,33,33,33},
							'{33,33,33,33,33,33,33,16,16,16,16,0,0,27,30,30,10,32,28,28,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,28,33,31,26,30,27,26,0,32,16,16,16,16,33,33,33,33,33},
							'{33,33,33,33,33,33,33,16,21,16,33,0,0,19,27,0,10,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,0,30,19,30,0,33,33,21,25,33,33,33,33,33,33},
							'{33,33,33,33,33,33,21,15,0,15,21,33,33,0,30,19,28,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,19,27,0,32,33,16,21,0,0,21,16,33,33,33,33},
							'{33,33,33,33,33,33,21,2,0,21,21,33,33,0,30,19,28,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,20,27,0,32,33,25,21,0,0,21,16,33,33,33,33},
							'{33,33,33,33,21,21,33,32,0,32,33,19,19,0,30,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,0,30,19,33,33,0,30,33,16,21,33,33,33},
							'{33,33,33,33,16,16,33,10,0,10,33,1,20,10,32,28,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,31,30,27,20,33,28,0,0,33,16,16,31,32,33},
							'{33,33,30,0,33,33,21,21,21,0,0,33,33,33,33,19,28,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,19,20,33,33,33,30,0,21,21,21,31,33,10,0,33},
							'{33,33,32,32,16,16,16,10,2,0,0,10,32,33,33,28,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,28,33,33,33,10,0,0,0,2,16,16,16,10,32,33},
							'{33,33,33,33,21,25,33,32,0,0,0,0,0,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,10,0,0,0,0,30,33,16,21,16,33,33},
							'{33,33,33,33,0,0,21,16,33,30,0,32,33,20,28,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,20,28,33,0,0,33,32,21,15,0,33,33,33},
							'{33,33,33,33,0,0,21,16,33,30,0,33,33,19,20,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,19,28,33,30,0,33,33,21,2,0,32,33,33},
							'{33,33,30,0,33,33,0,0,21,16,33,0,0,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,32,0,33,33,21,21,0,10,33,10,0,33},
							'{33,33,10,30,33,33,0,2,15,16,33,30,26,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,32,26,32,33,15,21,0,32,33,32,30,33},
							'{33,33,33,33,33,33,21,16,33,10,0,19,19,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,28,19,26,0,33,33,21,16,33,33,33,33},
							'{33,33,33,33,33,33,21,16,33,10,0,19,20,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,28,19,26,0,33,33,21,16,33,33,33,33},
							'{33,33,33,33,33,33,21,16,33,10,0,19,19,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,28,19,26,0,33,33,21,31,33,33,33,33},
							'{33,33,32,10,33,33,0,15,16,32,32,30,10,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,32,30,32,32,16,15,2,10,33,32,10,33},
							'{33,33,30,0,33,33,0,0,21,16,33,0,0,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,32,0,33,33,21,21,0,10,33,10,0,33},
							'{33,33,33,33,0,0,21,16,33,10,0,33,33,20,1,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,19,28,33,30,0,33,16,21,0,0,31,33,33},
							'{33,33,33,33,0,0,21,32,33,30,0,33,33,19,1,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,19,28,33,30,0,33,33,21,18,0,32,33,33},
							'{33,33,33,33,21,16,33,32,0,0,0,0,0,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,10,0,0,0,0,0,33,16,21,33,33,33},
							'{33,33,33,28,16,15,33,10,0,0,0,30,10,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,32,30,0,0,0,30,16,16,10,31,32,33},
							'{33,33,30,0,33,33,21,21,21,0,0,33,33,33,33,19,28,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,19,20,33,33,33,30,0,21,21,21,16,33,10,0,33},
							'{33,33,32,32,16,16,16,10,2,10,32,28,28,32,10,28,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,28,33,32,31,28,32,10,0,2,16,16,16,32,32,33},
							'{33,33,33,33,21,25,33,32,0,32,33,20,19,0,30,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,0,27,19,33,33,0,30,33,16,21,16,33,33},
							'{33,33,33,33,33,16,25,21,0,15,25,33,33,0,30,20,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,20,10,0,10,33,31,21,0,0,21,16,33,33,33,33},
							'{33,33,33,33,33,33,21,0,0,2,21,33,33,0,30,19,28,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,19,27,0,10,33,16,21,0,0,21,31,33,33,33,33},
							'{33,33,33,33,33,33,33,16,21,16,33,0,0,19,27,0,32,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,0,30,19,30,0,33,33,21,25,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,16,15,16,33,0,0,19,30,26,32,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,26,30,19,26,0,32,33,21,16,33,33,33,33,33,33},
							'{33,33,33,33,33,33,21,16,33,16,21,0,0,0,30,19,30,0,19,19,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,1,19,0,0,19,27,0,0,0,21,21,33,33,21,16,33,33,33,33},
							'{33,33,33,33,33,33,16,33,33,16,16,0,2,10,10,25,30,0,30,27,16,33,33,33,28,33,33,33,33,28,28,28,33,33,33,33,28,33,33,33,16,10,27,0,0,25,10,10,0,0,10,16,33,33,16,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,21,21,33,33,21,0,0,0,0,21,21,33,28,19,33,33,33,33,19,19,19,28,33,33,33,19,20,33,16,21,0,0,0,0,21,16,33,16,21,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,10,28,33,33,33,30,0,33,16,21,0,0,0,0,19,1,33,28,19,31,16,33,33,33,28,28,33,33,16,16,19,20,33,33,19,30,0,0,0,21,15,33,10,0,33,33,33,33,10,33,33,33,33,33},
							'{33,33,33,33,33,33,0,10,33,33,33,0,0,33,33,21,2,0,0,0,19,20,33,28,19,25,21,33,33,33,33,33,33,33,21,21,19,20,33,28,19,30,0,0,0,21,16,33,10,0,33,33,33,33,0,10,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,16,0,10,33,0,0,19,19,0,32,33,30,0,20,20,0,0,0,27,20,30,0,33,33,0,27,19,26,0,33,33,0,10,33,33,33,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,0,32,33,30,0,19,19,0,10,33,10,0,19,19,0,0,0,30,19,30,0,33,28,0,30,19,30,0,33,33,0,10,33,33,33,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,21,21,33,33,33,16,21,33,33,21,21,21,0,0,31,33,0,0,21,21,21,0,0,33,33,0,0,21,21,21,16,33,21,21,33,33,33,16,21,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,16,16,28,33,33,16,16,32,33,16,15,2,15,30,32,33,0,0,31,16,15,15,0,32,16,30,30,0,21,31,32,33,16,31,33,33,33,10,16,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,33,33,0,10,33,33,33,30,0,33,33,0,10,33,16,21,0,0,33,33,33,10,0,21,21,33,33,0,10,33,10,0,33,33,33,28,0,32,33,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,33,33,32,28,33,33,16,10,32,33,33,32,33,33,16,21,10,32,16,16,16,32,32,21,21,33,33,32,33,33,33,10,16,16,33,33,10,33,33,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,16,21,33,33,33,33,33,33,33,16,21,33,33,21,21,21,16,33,15,21,33,33,33,33,33,33,33,21,21,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,3,16,33,33,33,15,30,33,33,33,10,30,16,33,33,33,3,16,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,21,16,33,33,33,0,0,33,33,33,10,0,33,33,33,33,21,16,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
							'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33}};
	end
	
	always_ff @ (posedge vsync_slow[3]) begin
		// When enable goes on iterate through the explosion textures:
		if(enable1 == 0) released1 <= 0;
		if(enable1 == 1 && released1 == 0) begin
			counter1 <= 1;
			released1 <= 1;
		end
		if(counter1 != 0) counter1 <= counter1 + 1;
		if(counter1 >= 2) counter1 <= 0;
		
		// 
		if(enable2 == 0) released2 <= 0;
		if(enable2 == 1 && released2 == 0) begin
			counter2 <= 1;
			released2 <= 1;
		end
		if(counter2 != 0) counter2 <= counter2 + 1;
		if(counter2 >= 2) counter2 <= 0;
		
		//
		if(enable3 == 0) released3 <= 0;
		if(enable3 == 1 && released3 == 0) begin
			counter3 <= 1;
			released3 <= 1;
		end
		if(counter3 != 0) counter3 <= counter3 + 1;
		if(counter3 >= 2) counter3 <= 0;
	end
	
	always_comb begin
		// Defaults:
		color = 0;
		draw = 0;
		
		// Make sure that the pointer is inside the normal bullet:
		//Explosion Animation 1:
		if(vga_x >= exp1_x && vga_x < exp1_x + width1 && vga_y >= exp1_y && vga_y < exp1_y + height1 && counter1 == 1) begin
		   // If the color is not pink output draw:
			if(explosion1[vga_y - exp1_y][vga_x - exp1_x] != 8 && explosion1[vga_y - exp1_y][vga_x - exp1_x] != 33) begin
			    draw = 1'b1;
			    color = explosion1[vga_y - exp1_y][vga_x - exp1_x];
			end
		end
		if(vga_x >= exp1_x && vga_x < exp1_x + width2 && vga_y >= exp1_y && vga_y < exp1_y + height2 && counter1 == 2) begin
		   // If the color is not pink output draw:
			if(explosion2[vga_y - exp1_y][vga_x - exp1_x] != 8 && explosion2[vga_y - exp1_y][vga_x - exp1_x] != 33) begin
			    draw = 1'b1;
			    color = explosion2[vga_y - exp1_y][vga_x - exp1_x];
			end
		end
		
		// Explosion Animation 2:
		if(vga_x >= exp2_x && vga_x < exp2_x + width1 && vga_y >= exp2_y && vga_y < exp2_y + height1 && counter2 == 1) begin
		   // If the color is not pink output draw:
			if(explosion1[vga_y - exp2_y][vga_x - exp2_x] != 8 && explosion1[vga_y - exp2_y][vga_x - exp2_x] != 33) begin
			    draw = 1'b1;
			    color = explosion1[vga_y - exp2_y][vga_x - exp2_x];
			end
		end
		if(vga_x >= exp2_x && vga_x < exp2_x + width2 && vga_y >= exp2_y && vga_y < exp2_y + height2 && counter2 == 2) begin
		   // If the color is not pink output draw:
			if(explosion2[vga_y - exp2_y][vga_x - exp2_x] != 8 && explosion2[vga_y - exp2_y][vga_x - exp2_x] != 33) begin
			    draw = 1'b1;
			    color = explosion2[vga_y - exp2_y][vga_x - exp2_x];
			end
		end
		
		// Explosion Animation 3:
		if(vga_x >= exp3_x && vga_x < exp3_x + width1 && vga_y >= exp3_y && vga_y < exp3_y + height1 && counter3 == 1) begin
		   // If the color is not pink output draw:
			if(explosion1[vga_y - exp3_y][vga_x - exp3_x] != 8 && explosion1[vga_y - exp3_y][vga_x - exp3_x] != 33) begin
			    draw = 1'b1;
			    color = explosion1[vga_y - exp3_y][vga_x - exp3_x];
			end
		end
		if(vga_x >= exp3_x && vga_x < exp3_x + width2 && vga_y >= exp3_y && vga_y < exp3_y + height2 && counter3 == 2) begin
		   // If the color is not pink output draw:
			if(explosion2[vga_y - exp3_y][vga_x - exp3_x] != 8 && explosion2[vga_y - exp3_y][vga_x - exp3_x] != 33) begin
			    draw = 1'b1;
			    color = explosion2[vga_y - exp3_y][vga_x - exp3_x];
			end
		end
	end
endmodule