library verilog;
use verilog.vl_types.all;
entity testbench_8 is
end testbench_8;
