//--------------------------------------------------------------------------------------------
// Sprite Mapper:
//
//		The sprite mapper is a glorified color mapper and it will draw the sprites with the 
//		top left corner at the (x,y) coordinate. The background moves based on the position of
//		samus. (She is in the middle on the screen)
//
//--------------------------------------------------------------------------------------------
// Pallate: (0,0,0), (0,0,255), (102,102,102), (0,255,255),(0,255,0), (64,128,0),(255,0,0),(255,102,102),(128,0,0),(248,146,56),(232,146,41),(27,175,0),(19,137,13),(255,49,62),(234,228,94),(126,0,246),(47,151,209),(156,89,33),(82,105,250),(43,93,83),(13,65,63),(37,75,258),(148,148,118),(60,70,17),(63,71,73),(34,28,28),(4,35,248),(186,0,37),(126,0,246),(103,0,183)
module sprite_mapper(
input logic clk, reset,
input logic [9:0] vgaX, vgaY, 
output logic [7:0] red, green, blue
);

	// Internal Signals:
	logic [6:0] bg_color;
	logic [6:0] powerUp_color;
	logic [6:0] bullet_color;
	logic [6:0] monster_color;
	logic [6:0] samus_color;
   logic [6:0] color;
	logic bulletDraw, monsterDraw, samusDraw, powerUpDraw;
	logic tempFlash;
	
	always_ff @(posedge clk) begin
	    if(vgaY == 479 && vgaX == 639) tempFlash <= ~tempFlash;
	end
 
	// This module acts as a mux on all of the different levels of sprites:

   // Texture Units:
	background bg(.background_start_addr(1'b0), .vga_x(vgaX), .vga_y(vgaY), .color(bg_color));
   bullet bull(.enable1(flash), .enable2(flash), .enable3(flash), 
		.vga_x(vgaX), .vga_y(vgaY), 
		.sprite1_x(120), .sprite1_y(40), 
		.sprite2_x(80), .sprite2_y(40), 
		.sprite3_x(40), .sprite3_y(40), 
		.sprite_num(1'b0),
		.color(bullet_color),
		.draw(bulletDraw));
	
	
	// Select the color based on priority:
	always_comb begin
	   // Default:
	   color = bg_color;	
		
		if(bulletDraw == 1'b1) color = bullet_color;
		else color = bg_color;
	end
	
	// Pass the color to pallate to output the proper color:
	always_comb begin
		//Defaults:
		red = 8'b0;
		green = 8'b0;
		blue = 8'b0;
		
		case(color)
			//Color 1:
			1: begin
				red = 44;
				green = 92;
				blue = 10;
			end
			//Color 2:
			2: begin
			//248,146,56
				red = 248;
				green = 146;
				blue = 56;
			end
			//Color 3:
			3: begin
			//(156,0,18
				red = 156;
				green = 0;
				blue = 18;
			end
			//Color 4:
			4: begin
			// 0, 255, 128
				red = 0;
				green = 255;
				blue = 128;
			end
			//Color 5:
			5: begin
			// 0,0,128
				red = 0;
				green = 0;
				blue = 128;
			end
			//Color 6:
			6: begin
			// 0,128,255
				red = 0;
				green = 128;
				blue = 255;
			end
			//Color 7:
			7: begin
			// 255,255,255
				red = 255;
				green = 255;
				blue = 255;
			end
			//Color 8:
			8: begin
				red = 0;
				green = 0;
				blue = 0;
			end
			//Color 9:
			9: begin
				red = 0;
				green = 0;
				blue = 255;
			end
			//Color 10:
			10: begin
				red = 102;
				green = 102;
				blue = 102;
			end
			//Color 11:
			11: begin
				red = 0;
				green = 255;
				blue = 255;
			end
			//Color 12
			12: begin
				red = 0;
				green = 255;
				blue = 0;
			end
			//Color 13:
			13: begin
				red = 64;
				green = 128;
				blue = 0;
			end
			//Color 14:
			14: begin
				red = 255;
				green = 0;
				blue = 0;
			end
			//Color 15:
			15: begin
				red = 255;
				green = 102;
				blue = 102;
			end
			//Color 16
			16: begin
				red = 128;
				green = 0;
				blue = 0;
			end
			//Color 17:
			17: begin
				red = 248;
				green = 146;
				blue = 56;
			end
			//Color 18:
			18: begin
				red = 232;
				green = 146;
				blue = 41;
			end
			//Color 19:
			19: begin
				red = 27;
				green = 175;
				blue = 0;
			end
			//Color 20:
			20: begin
				red = 19;
				green = 137;
				blue = 13;
			end
			//Color 21:
			21: begin
				red = 255;
				green = 49;
				blue = 62;
			end
			//Color 22:
			22: begin
				red = 234;
				green = 228;
				blue = 94;
			end
			//Color 23:
			23: begin
				red = 126;
				green = 0;
				blue = 246;
			end
			//Color 24:
			24: begin
				red = 47;
				green = 151;
				blue = 209;
			end
			//Color 25:
			25: begin
				red = 156;
				green = 89;
				blue = 33;
			end
			//Color 26:
			26: begin
				red = 82;
				green = 105;
				blue = 250;
			end
			//Color 27:
			27: begin
				red = 43;
				green = 93;
				blue = 83;
			end
			//Color 28:
			28: begin
				red = 13;
				green = 65;
				blue = 63;
			end
			//Color 29:
			29: begin
				red = 37;
				green = 75;
				blue = 258;
			end
			//Color 30:
			30: begin
				red = 148;
				green = 148;
				blue = 118;
			end
			//Color 31:
			31: begin
				red = 60;
				green = 70;
				blue = 17;
			end
			//Color 32:
			32: begin
				red = 63;
				green = 71;
				blue = 73;
			end
			//Color 33:
			33: begin
				red = 34;
				green = 28;
				blue = 28;
			end
			34: begin
				red = 4;
				green = 35;
				blue = 248;
			end
			35: begin
				red = 186;
				green = 0;
				blue = 37;
			end
			36: begin
				red = 103;
				green = 0;
				blue = 246;
			end
			37: begin
				red = 103;
				green = 0;
				blue = 183;
			end
			// Default:
			default: begin
				red = 0;
				green = 0;
				blue = 0;
			end
		endcase
	end
	
endmodule

/*
//--------------------------------------------------------------------------------------------
// Samus:
//
//		If the vga pixel pointer is within the samus sprite, return a proper color:
//		Priority 1
//
//--------------------------------------------------------------------------------------------
module samus(
	input logic  			enable,
	input logic  [10:0] 	vga_x, vga_y, sprite_x, sprite_y,
	input logic  [1:0] 	sprite_num,
	output logic [5:0] 	color,
	output logic 			draw
);
	// Samus Sprites:
	parameter [9:0] height = 70;
	parameter [9:0] width = 45;
	
	// Samus Combinational Logic:
	always_comb begin
	   // Determine the width and height of the 
	   case(sprite_num)
		// SAMUS STAND:
		2b'00: begin
			// Output the "draw" signal:
			// Make sure that the pointer is inside the sprite:
			if(vga_x > sprite_x && vga_x < sprite_x + width && vga_y > sprite_y && vga_y < sprite_y + height) begin
				// If the color is not pink output draw:
				//if( != 63)
				draw = 1'b1;
				color = 6'b0;
			end
			else begin
				draw = 1'b0;
				color = 6'b0;
			end
		end
		// SAMUS WALK 1:
		2'b01: begin
			// Output the "draw" signal:
			// Make sure that the pointer is inside the sprite:
			if(vga_x > sprite_x && vga_x < sprite_x + width && vga_y > sprite_y && vga_y < sprite_y + height) begin
				// If the color is not pink output draw:
				//if( != 63)
				draw = 1'b1;
				color = 6'b0;
			end
			else begin
				draw = 1'b0;
				color = 6'b0;
			end
		end
		// SAMUS WALK 2:
		2'b10: begin
			// Output the "draw" signal:
			// Make sure that the pointer is inside the sprite:
			if(vga_x > sprite_x && vga_x < sprite_x + width && vga_y > sprite_y && vga_y < sprite_y + height) begin
				// If the color is not pink output draw:
				//if( != 63)
				draw = 1'b1;
				color = 6'b0;
			end
			else begin
				draw = 1'b0;
				color = 6'b0;
			end
		end
		// SAMUS WALK 3:
		2'b11: begin
			// Output the "draw" signal:
			// Make sure that the pointer is inside the sprite:
			if(vga_x > sprite_x && vga_x < sprite_x + width && vga_y > sprite_y && vga_y < sprite_y + height) begin
				// If the color is not pink output draw:
				//if( != 63)
				draw = 1'b1;
				color = 6'b0;
			end
			else begin
				draw = 1'b0;
				color = 6'b0;
			end
		end
		endcase
	end
endmodule


//--------------------------------------------------------------------------------------------
// Monster:
//
//		If the vga pixel pointer is within the monster(s), return a proper color:
//		Priority 2
//		
//--------------------------------------------------------------------------------------------
module monster(
	input logic  			enable1, enable2, enable3,
	input logic  [10:0] 	vga_x, vga_y, sprite1_x, sprite1_y, sprite2_x, sprite2_y, sprite3_x, sprite3_y,
	input logic  [1:0] 	sprite_num,
	output logic [5:0] 	color,
	output logic 			draw
);
	// Monster Sprites:
	parameter [9:0] height = 70;
	parameter [9:0] width = 45;
	
	// Monster Combinational Logic:
	always_comb begin
		// Make sure that the pointer is inside the MONSTER 1:
		if(vga_x > sprite1_x && vga_x < sprite1_x + width && vga_y > sprite1_y && vga_y < sprite1_y + height && enable1) begin
		   // If the color is not pink output draw:
			//if( != 63)
			draw = 1'b1;
			color = 6'b0;
		end
		else begin
			draw = 1'b0;
			color = 6'b0;
		end
		// MONSTER 2
		if(vga_x > sprite2_x && vga_x < sprite2_x + width && vga_y > sprite2_y && vga_y < sprite2_y + height && enable2) begin
		   // If the color is not pink output draw:
			//if( != 63)
			draw = 1'b1;
			color = 6'b0;
		end
		else begin
			draw = 1'b0;
			color = 6'b0;
		end
		// MONSTER 3
		if(vga_x > sprite1_x && vga_x < sprite1_x + width && vga_y > sprite1_y && vga_y < sprite1_y + height && enable3) begin
		   // If the color is not pink output draw:
			//if( != 63)
			draw = 1'b1;
			// Chose the proper color:
			color = 6'b0;
		end
		else begin
			draw = 1'b0;
			color = 6'b0;
		end
	end
endmodule


//--------------------------------------------------------------------------------------------
// PowerUp:
//
//		If the vga pixel pointer is within the powerUp, return a proper color:
//		Priority 3
//		
//--------------------------------------------------------------------------------------------
module power_up(
	input logic  			enable1, enable2, enable3,
	input logic  [10:0] 	vga_x, vga_y, sprite1_x, sprite1_y, sprite2_x, sprite2_y, sprite3_x, sprite3_y,
	input logic  [1:0] 	sprite_num,
	output logic [5:0] 	color,
	output logic 			draw
);
// Mux the certain power up:
// powerUp Sprites:
	parameter [9:0] height = 70;
	parameter [9:0] width = 45;
	
	// Monster Combinational Logic:
	always_comb begin
		// Make sure that the pointer is inside the powerUp 1:
		if(vga_x > sprite1_x && vga_x < sprite1_x + width && vga_y > sprite1_y && vga_y < sprite1_y + height && enable1) begin
		   // If the color is not pink output draw:
			//if( != 63)
			draw = 1'b1;
			color = 6'b0;
		end
		else begin
			draw = 1'b0;
			color = 6'b0;
		end
		// powerUp 2
		if(vga_x > sprite2_x && vga_x < sprite2_x + width && vga_y > sprite2_y && vga_y < sprite2_y + height && enable2) begin
		   // If the color is not pink output draw:
			//if( != 63)
			draw = 1'b1;
			color = 6'b0;
		end
		else begin
			draw = 1'b0;
			color = 6'b0;
		end
		// powerUp 3
		if(vga_x > sprite1_x && vga_x < sprite1_x + width && vga_y > sprite1_y && vga_y < sprite1_y + height && enable3) begin
		   // If the color is not pink output draw:
			//if( != 63)
			draw = 1'b1;
			// Chose the proper color:
			color = 6'b0;
		end
		else begin
			draw = 1'b0;
			color = 6'b0;
		end
	end
endmodule
*/

//--------------------------------------------------------------------------------------------
// Bullet:
//
//		If the vga pixel pointer is within the bullet(s), return a proper color:
//		Priority 4
//		
//--------------------------------------------------------------------------------------------
module bullet(
	input logic  			enable1, enable2, enable3,
	input logic  [10:0] 	vga_x, vga_y, sprite1_x, sprite1_y, sprite2_x, sprite2_y, sprite3_x, sprite3_y,
	input logic  [1:0] 	sprite_num,
	output logic [5:0] 	color,
	output logic 			draw
);
// Mux the bullet instances:
// powerUp Sprites:
	parameter [9:0] height = 10;
	parameter [9:0] width = 10;
	
	int BulletN [10][10];
	int BulletE [10][10];
	
	always_ff begin
	    BulletN = '{'{00,00,00,00,06,06,00,00,00,00},
		             '{00,00,06,06,06,06,06,06,00,00},
						 '{00,06,06,06,06,06,06,06,06,00},
						 '{00,06,06,06,06,06,06,06,06,00},
						 '{06,06,06,06,06,06,06,06,06,06},
						 '{06,06,06,06,06,06,06,06,06,06},
						 '{00,06,06,06,06,06,06,06,06,00},
						 '{00,06,06,06,06,06,06,06,06,00},
						 '{00,00,06,06,06,06,06,06,00,00},
						 '{00,00,00,00,06,06,00,00,00,00}};
		/* BulletE = '{'{63,63,63,63,06,06,63,63,63,63},
		             '{63,63,06,06,06,06,06,06,63,63},
						 '{63,06,06,06,06,06,63,63,06,63},
						 '{63,06,06,06,06,06,63,63,06,63},
						 '{06,06,06,06,06,06,63,63,63,06},
						 '{06,06,06,06,06,06,63,63,63,06},
						 '{63,06,06,06,06,06,63,63,63,63},
						 '{63,06,63,06,06,06,63,63,63,63},
						 '{63,63,06,06,06,06,63,63,63,63},
						 '{63,63,63,63,06,06,63,63,63,63}}; */
	end
	
	// Monster Combinational Logic:
	always_comb begin
	// Defaults:
	color = 0;
	draw = 0;
		// Make sure that the pointer is inside the normal bullet:
		if(vga_x > sprite1_x && vga_x < sprite1_x + width && vga_y > sprite1_y && vga_y < sprite1_y + height && enable1) begin
		   // If the color is not pink output draw:
			if(BulletN[vga_x - sprite1_x][vga_y - sprite1_y] != 0) begin
			    draw = 1'b1;
			    color = BulletN[vga_x - sprite1_x][vga_y - sprite1_y];
			end
		end
		else begin
			draw = 1'b0;
			color = 6'b0;
		end
		// powerUp 2
		if(vga_x > sprite2_x && vga_x < sprite2_x + width && vga_y > sprite2_y && vga_y < sprite2_y + height && enable2) begin
		   // If the color is not pink output draw:
			if(BulletN[vga_x - sprite2_x][vga_y - sprite2_y] != 0) begin
			    draw = 1'b1;
			    color = BulletN[vga_x - sprite2_x][vga_y - sprite2_y];
			end
		end
		else begin
			draw = 1'b0;
			color = 6'b0;
		end
		// powerUp 3
		if(vga_x > sprite3_x && vga_x < sprite3_x + width && vga_y > sprite3_y && vga_y < sprite3_y + height && enable3) begin
		   // If the color is not pink output draw:
			if(BulletN[vga_x - sprite3_x][vga_y - sprite3_y] != 0) begin
			    draw = 1'b1;
			    color = BulletN[vga_x - sprite3_x][vga_y - sprite3_y];
			end
		end
		else begin
			draw = 1'b0;
			color = 6'b0;
		end
	end
endmodule


//--------------------------------------------------------------------------------------------
// Background:
//
//		If the vga pixel pointer is within the proper background tile, return a proper color:
//		Priority 5
//		
//--------------------------------------------------------------------------------------------
module background(
   input logic  [10:0]	background_start_addr,
	input logic  [9:0] 	vga_x, vga_y,
	output logic [5:0] 	color
);
	// Background Tile sizes:
	parameter [9:0] height = 30;
	parameter [9:0] width = 30;
	parameter [9:0] screenH = 16;
	parameter [9:0] screenW = 22;
	// Combinational math an returns 
	logic [10:0] background_x, background_y; // Normalized background array pointers:
	logic [10:0] tile_x, tile_y; // Normalized tile coordinate pointers:
	
	// Sprites: 8 different backgrounds:
	int BG1 [height][width];
	int BG2 [height][width];
	int BG3 [height][width];
	int BG4 [height][width];
	int BG5 [height][width];
	int BG6 [height][width];
	int BG7 [height][width];
	int BG8 [height][width];
	int dummy [screenH][screenW];
	
	//-------------------------------------------------------------------------------------------------------------
	// Sprite arrays + dummy background array:
	//-------------------------------------------------------------------------------------------------------------
	always_ff begin
		dummy = '{'{1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1},
		          '{1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1},
					 '{1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1},
					 '{1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1},
					 '{1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,4,4,4,0,1,1},
					 '{1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,5,5,5,0,1,1},
					 '{1,0,0,0,0,0,0,1,2,3,3,0,0,0,0,0,6,6,6,0,1,1},
					 '{1,0,0,0,0,0,0,3,2,2,2,0,0,0,0,0,7,7,7,0,1,1},
					 '{1,0,0,0,0,1,1,1,1,0,3,0,0,0,0,0,0,0,0,0,1,1},
					 '{1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1},
					 '{1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1},
					 '{1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1},
					 '{1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1},
					 '{1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1},
					 '{1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1},
					 '{1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1}};
		// All Black (08):
		BG1 = '{'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
		        '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33}};
		// BLue_brick1:
		BG2 = '{'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
		        '{33,33,33,33,33,33,33,28,33,28,33,28,33,28,33,28,33,28,33,28,33,28,33,28,33,28,33,33,33,33},
				  '{33,33,33,33,33,28,24,26,24,26,24,26,24,26,24,26,24,26,24,26,24,26,24,26,24,26,26,33,33,33},
				  '{33,33,28,28,28,29,29,29,29,29,29,29,29,29,29,29,29,29,29,29,29,29,29,29,29,29,29,33,33,33},
				  '{33,33,26,24,26,26,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,33,33,33},
				  '{33,33,26,26,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,33,33,33},
				  '{33,33,26,26,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,33,33,33},
				  '{33,33,26,26,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,33,33,33},
				  '{33,33,26,26,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,05,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,28,28,28,28,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,28,24,26,24,26,26,33,33,33},
				  '{33,33,28,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,33,33,33,28,26,26,29,29,34,33,33,33},
              '{33,33,26,24,26,24,26,24,26,24,26,24,26,24,26,24,26,26,33,33,33,28,24,29,34,34,34,33,33,33},
              '{33,33,26,26,29,34,29,34,34,29,34,34,29,34,34,29,34,34,33,33,26,29,34,34,34,34,34,33,33,33},
				  '{33,33,26,26,34,34,34,34,34,34,34,34,34,34,34,34,34,34,33,33,26,26,34,34,34,34,34,33,33,33},
				  '{33,33,26,26,34,34,34,34,34,34,34,34,34,34,34,34,34,34,33,33,24,29,34,34,34,34,34,33,33,33},
				  '{33,33,26,26,34,34,34,34,34,34,34,34,34,34,34,34,5,5,33,33,26,26,34,34,34,34,34,33,33,33},
				  '{33,33,26,26,34,34,34,34,34,34,34,34,34,34,34,34,33,33,33,33,26,26,34,34,34,34,34,33,33,33},
				  '{33,33,28,28,5,33,5,33,5,33,5,33,5,33,5,33,33,33,33,33,28,34,33,5,33,5,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,26,26,26,26,26,26,26,33,33,33,33,33,33,33,33,33,33,33,26,26,26,26,26,26,27,33,33,33},
				  '{33,33,26,24,26,24,26,24,26,33,33,33,33,33,33,33,33,33,33,33,26,24,26,24,26,24,26,33,33,33},
				  '{33,33,26,26,34,34,34,34,34,34,34,34,34,34,34,34,34,34,26,26,34,34,34,34,34,34,34,33,33,33},
				  '{33,33,26,26,34,34,34,34,34,34,34,34,34,34,34,34,34,34,26,26,34,34,34,34,34,34,34,33,33,33},
				  '{33,33,26,26,34,34,34,34,34,34,34,34,34,34,34,34,34,34,24,26,34,34,34,34,34,34,34,33,33,33},
				  '{33,33,28,27,5,5,5,5,5,5,5,5,5,5,5,5,5,5,27,28,5,5,5,5,5,5,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
				  '{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33}};
		
		// Brick grey:
		BG3 =     '{'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,33,33},
						'{33,33,33,33,33,33,10,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,26,33,33},
						'{33,33,33,26,26,26,22,26,30,26,22,30,26,22,30,26,22,30,26,22,30,26,22,30,26,22,30,10,33,33},
						'{33,33,33,7,7,7,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,10,33,33},
						'{33,33,33,7,22,30,30,30,30,30,10,30,30,10,30,30,10,30,30,10,30,30,10,30,30,10,30,10,33,33},
						'{33,33,33,7,7,10,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,10,33,33},
						'{33,33,33,7,7,10,30,30,30,10,30,10,30,30,10,30,30,10,30,30,10,30,30,10,30,30,30,10,33,33},
						'{33,33,33,10,10,32,32,31,32,32,31,10,31,32,31,32,31,32,31,32,31,32,31,32,31,32,31,31,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,32,30,30,30,30,10,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,10,7,7,7,7,26,33,33},
						'{33,33,33,26,22,26,7,26,22,26,7,26,22,26,7,26,22,26,22,33,33,33,10,7,26,30,30,10,33,33},
						'{33,33,33,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,26,33,33,33,10,7,30,30,30,10,33,33},
						'{33,33,33,7,7,10,30,30,10,30,30,10,30,30,10,30,30,30,10,33,31,7,26,30,30,30,30,10,33,33},
						'{33,33,33,7,22,30,30,30,30,30,30,30,30,30,30,30,10,30,10,33,32,7,22,30,30,30,30,10,33,33},
						'{33,33,33,7,7,10,30,30,30,10,30,10,30,10,30,30,30,30,10,33,32,7,26,30,30,10,30,10,33,33},
						'{33,33,33,7,26,30,30,30,30,30,30,30,30,30,10,30,10,31,33,33,32,7,22,30,30,30,30,10,33,33},
						'{33,33,33,7,7,10,30,10,30,10,30,30,10,30,30,30,30,33,33,33,32,7,26,30,30,30,30,10,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,7,7,7,7,7,7,7,33,33,33,33,33,33,33,33,33,33,31,7,7,7,7,7,7,26,33,33},
						'{33,33,33,7,7,7,7,7,7,26,33,33,33,33,33,33,33,33,33,33,10,7,7,7,7,7,22,26,33,33},
						'{33,33,33,7,7,10,10,30,30,30,30,30,30,30,30,30,30,30,30,7,7,10,10,10,10,10,30,10,33,33},
						'{33,33,33,7,22,10,30,30,30,30,30,30,30,30,30,30,30,30,30,7,26,30,30,30,30,30,30,10,33,33},
						'{33,33,33,7,7,10,30,30,30,30,30,30,10,30,10,30,10,30,30,7,22,30,30,30,30,10,30,10,33,33},
						'{33,33,33,32,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,32,32,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33}};
		// Brick green:
		BG4 =     '{'{33,33,33,32,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,32,32,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,31,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,33,33,33},
						'{33,33,33,33,33,31,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,25,33,33,33},
						'{33,33,18,18,18,13,20,19,19,20,19,19,19,19,19,19,19,19,19,20,19,19,19,19,20,19,20,33,33,33},
						'{33,33,18,18,25,27,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,33,33,33},
						'{33,33,18,18,19,20,20,19,20,19,20,19,20,19,20,19,20,20,19,20,19,20,20,19,20,20,20,33,33,33},
						'{33,33,18,18,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,19,20,20,19,20,20,33,33,33},
						'{33,33,18,18,19,20,20,19,20,19,20,19,20,19,20,20,20,19,20,19,20,20,20,19,20,20,20,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,31,18,18,18,18,18,33,33,33},
						'{33,33,33,16,33,31,33,16,33,31,33,16,33,31,33,16,33,31,33,33,33,31,18,18,13,18,25,33,33,33},
						'{33,33,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,33,33,33,31,18,19,20,20,20,33,33,33},
						'{33,33,18,18,13,27,25,13,27,25,13,27,25,27,13,25,27,25,33,33,31,25,25,19,20,19,20,33,33,33},
						'{33,33,18,18,20,20,20,20,20,20,20,20,19,20,20,20,19,20,33,33,18,13,20,20,20,20,20,33,33,33},
						'{33,33,18,18,19,20,19,20,19,20,19,20,20,20,19,20,20,20,33,33,18,25,19,20,19,20,20,33,33,33},
						'{33,33,18,18,19,20,20,20,20,20,20,20,20,20,20,19,20,20,33,33,18,13,20,20,20,20,20,33,33,33},
						'{33,33,18,18,19,20,19,20,19,20,20,20,19,20,20,20,33,33,33,33,18,25,19,20,19,20,20,33,33,33},
						'{33,33,25,25,20,28,20,27,20,27,20,27,20,27,20,20,33,33,33,33,18,31,20,28,20,28,28,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,31,31,31,31,31,31,31,33,33,33,33,33,33,33,33,33,33,33,31,31,31,31,31,31,31,33,33,33},
						'{33,33,18,18,18,18,18,18,18,33,33,33,33,33,33,33,33,33,33,33,18,18,18,18,18,18,18,33,33,33},
						'{33,33,18,18,19,27,19,27,19,28,28,28,28,28,28,28,28,28,25,25,27,19,27,19,27,19,27,33,33,33},
						'{33,33,18,18,19,20,20,20,20,19,20,19,19,20,19,19,20,19,18,18,20,20,20,20,20,20,20,33,33,33},
						'{33,33,18,18,20,20,19,20,20,20,20,20,20,20,20,20,20,20,18,18,19,20,20,19,20,20,20,33,33,33},
						'{33,33,18,25,20,20,20,20,20,20,20,20,20,20,20,20,20,20,18,25,20,20,20,20,20,20,28,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33},
						'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33}};
		// Blue door bot mid 1:
		BG5 =     '{'{3,34,29,29,34,29,34,29,34,29,34,29,34,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{2,29,29,29,29,29,29,29,29,29,29,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{25,29,34,29,29,34,29,29,34,29,29,29,34,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,34,29,29,29,29,29,29,29,29,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,29,34,29,34,29,34,29,29,29,29,29,29,34,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,34,29,29,29,29,29,29,34,29,34,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,29,34,29,29,29,34,29,29,29,29,29,34,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,34,29,29,34,29,29,29,29,34,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,29,34,29,29,29,29,34,29,29,29,34,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,34,29,29,29,34,29,29,29,29,29,29,29,34,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,29,34,29,29,29,29,29,34,29,29,34,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,34,29,29,29,34,29,29,29,29,29,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,29,34,29,29,29,29,34,29,34,29,34,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,34,29,29,34,29,29,29,29,29,29,29,29,34,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,29,34,29,29,29,34,29,29,34,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{18,29,29,29,29,29,29,29,29,29,29,34,29,34,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{18,29,34,29,34,29,29,34,29,34,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,34,29,29,29,29,29,29,29,29,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,29,34,29,29,34,29,34,29,29,34,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,29,29,29,29,29,29,29,29,29,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,29,34,29,29,34,29,29,34,29,34,29,34,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,29,29,29,29,29,29,29,29,29,29,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{3,34,29,29,34,29,34,29,34,29,29,34,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,34,29,29,29,29,29,29,29,29,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{3,34,29,34,29,29,34,29,29,34,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,34,29,29,29,29,29,29,29,29,29,34,29,34,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{3,34,29,29,34,29,29,34,29,34,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,34,29,29,29,29,29,29,29,29,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{16,34,29,29,34,29,34,29,29,34,29,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
						'{21,29,29,29,29,29,29,29,29,29,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}};
		// Blue Door Bot Right:
		BG6 =  '{'{21,29,29,29,29,29,29,29,29,29,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{2,29,34,29,29,34,29,34,29,34,29,29,29,34,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,29,29,29,29,29,29,29,29,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,29,34,29,29,34,29,29,34,29,34,29,34,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,29,29,29,29,29,29,29,29,29,28,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,34,29,34,29,34,29,29,34,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,34,29,29,29,29,29,29,29,29,29,29,5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,29,34,29,29,34,29,29,34,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,34,29,29,29,29,29,29,29,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,34,29,34,29,24,26,29,34,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,34,29,29,29,29,29,26,7,29,29,29,5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,29,29,34,29,26,7,34,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,34,29,29,29,29,24,26,26,29,29,34,28,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,34,29,24,7,26,29,29,29,29,5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,29,29,29,29,24,7,29,29,34,29,34,33,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{2,29,29,34,29,34,24,7,26,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,29,29,26,26,7,7,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,34,24,7,7,7,26,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,7,7,7,24,29,29,34,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,29,7,7,7,26,29,29,29,34,28,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,7,7,7,24,34,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,29,7,7,26,26,29,34,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,7,26,34,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,29,24,26,29,29,34,28,5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,34,29,34,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,34,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,28,34,28,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}};
		// Blue Door bottop:
		BG7 =  '{'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{31,28,5,5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{2,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,34,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,34,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,29,29,34,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,29,29,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,7,26,29,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,29,7,26,24,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,7,7,7,24,29,34,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,29,7,7,7,26,29,29,34,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,7,7,7,24,29,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,29,29,24,7,7,7,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,26,7,7,7,26,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,34,29,34,29,24,7,26,34,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,29,29,29,34,24,7,26,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{2,29,34,29,29,29,24,7,29,29,29,34,29,5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{25,34,29,29,34,29,26,26,24,24,34,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,29,29,29,29,26,7,29,29,29,5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,34,29,29,34,29,29,26,7,29,34,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,29,29,29,29,26,7,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,34,29,29,34,29,29,29,34,29,29,34,28,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,29,29,34,29,29,29,29,29,34,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,34,29,34,29,29,29,34,29,34,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,29,29,29,29,29,29,29,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,34,29,29,34,29,34,29,29,34,29,34,28,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,34,29,29,29,29,29,29,29,29,29,29,29,34,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,34,29,29,34,29,29,34,29,29,34,29,29,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{16,29,29,29,29,29,29,29,29,29,29,29,29,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{3,34,29,29,34,29,34,29,34,29,34,29,34,29,29,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}};
		// Blue Door left:
		BG8 =  '{'{33,21,21,21,25,21,21,25,21,21,25,21,21,21,21,21,21,21,21,25,21,21,25,21,21,21,25,21,21,29},
					'{16,18,2,2,2,2,2,2,2,2,2,2,2,18,2,18,2,18,2,2,2,2,2,2,2,2,2,2,2,29},
					'{33,2,10,29,24,29,24,29,29,24,29,24,29,16,16,2,30,29,24,29,29,24,29,24,29,29,24,32,16,29},
					'{16,2,24,29,29,29,29,29,29,29,29,29,24,16,16,2,30,29,29,29,29,29,29,29,29,24,29,33,16,29},
					'{33,2,10,29,33,16,16,16,16,16,16,28,29,16,16,18,30,29,28,16,16,16,16,16,16,28,29,28,16,34},
					'{16,2,24,29,16,16,32,33,32,16,16,26,29,16,16,2,30,29,28,16,16,28,32,16,16,10,24,33,16,34},
					'{33,2,24,29,33,16,29,29,24,26,2,24,29,16,16,2,30,29,28,16,29,29,29,24,2,10,29,28,16,29},
					'{16,2,10,29,16,16,29,24,29,24,2,24,29,16,16,2,10,29,28,16,29,24,29,24,18,10,29,31,16,34},
					'{33,2,24,29,33,16,29,29,24,26,2,24,29,16,16,2,30,29,28,16,28,29,29,24,18,10,24,28,16,29},
					'{16,2,24,29,16,16,30,30,30,18,2,26,29,16,16,2,30,29,28,16,25,30,30,18,2,26,29,28,16,34},
					'{33,2,10,29,28,16,2,18,2,2,2,24,29,16,16,2,10,29,28,16,2,2,2,2,2,10,29,28,16,29},
					'{16,2,24,29,29,24,29,29,29,24,29,29,24,16,16,2,30,29,24,29,29,29,29,24,29,24,29,28,16,34},
					'{33,18,10,29,29,28,29,29,29,28,29,29,29,16,16,18,25,29,29,29,29,27,29,29,29,34,29,16,16,29},
					'{33,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,34},
					'{33,21,16,25,16,25,16,25,16,25,16,25,3,25,21,16,25,3,25,16,25,16,25,3,25,16,25,21,16,29},
					'{33,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,18,2,2,29},
					'{16,2,10,26,26,24,26,24,26,24,26,24,26,25,16,2,18,24,26,24,26,24,26,24,26,24,24,10,16,29},
					'{33,2,10,29,24,29,29,29,24,29,29,29,24,16,3,2,30,29,29,24,29,29,29,24,29,29,29,31,16,34},
					'{16,2,24,29,28,16,16,16,16,33,16,29,29,16,16,18,30,29,28,16,33,16,16,16,33,28,29,28,16,34},
					'{33,2,24,29,16,16,16,16,16,16,16,28,29,16,16,2,30,29,28,16,16,16,16,16,3,32,29,31,16,29},
					'{16,2,10,29,33,16,29,29,24,26,2,24,29,16,16,2,10,29,28,16,29,29,29,24,18,10,24,28,16,34},
					'{33,2,24,29,16,16,24,29,29,24,2,26,29,16,16,2,30,29,28,16,29,24,29,24,2,26,29,28,16,29},
					'{16,2,24,29,28,16,29,24,29,24,2,24,29,16,16,2,30,29,28,16,28,29,24,29,2,10,29,28,16,34},
					'{33,2,10,29,16,16,10,26,10,30,18,24,29,16,16,2,10,29,28,16,10,10,26,10,2,10,24,28,16,29},
					'{16,2,24,29,33,16,2,2,2,2,2,26,29,16,16,2,30,29,28,16,21,2,2,2,2,10,29,28,16,34},
					'{33,2,24,29,29,29,26,24,26,26,24,29,24,16,16,18,30,29,29,29,26,24,26,24,29,24,29,28,16,29},
					'{16,2,10,29,24,29,29,29,24,29,29,24,29,16,16,2,10,24,29,24,29,29,29,24,29,29,24,33,16,34},
					'{33,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,29},
					'{33,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,34},
					'{33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33}};
	end
	
	
	always_comb begin
		// Determines the upper left corner of the tile sprite:
		// Defaults:
		background_x = 0;
		background_y = 0;
		tile_x = 0;
		tile_y = 0;
		
		if(vga_x >= 0 && vga_x < width) begin
	   	background_x = 0;
			tile_x = 0;
		end
		if(vga_x >= width && vga_x < 2*width) begin
			background_x = width;
			tile_x = 1;
		end
		if(vga_x >= 2*width && vga_x < 3*width) begin
			background_x = 2*width;
			tile_x = 2;
		end
		if(vga_x >= 3*width && vga_x < 4*width) begin
			background_x = 3*width;
			tile_x = 3;
		end
		if(vga_x >= 4*width && vga_x < 5*width) begin 
			background_x = 4*width;
			tile_x = 4;
		end
		if(vga_x >= 5*width && vga_x < 6*width) begin
			background_x = 5*width;
			tile_x = 5;
		end
		if(vga_x >= 6*width && vga_x < 7*width) begin
			background_x = 6*width;
			tile_x = 6;
		end
		if(vga_x >= 7*width && vga_x < 8*width) begin
			background_x = 7*width;
			tile_x = 7;
		end
		if(vga_x >= 8*width && vga_x < 9*width) begin
			background_x = 8*width;
			tile_x = 8;
		end
		if(vga_x >= 9*width && vga_x < 10*width) begin
			background_x = 9*width;
			tile_x = 9;
		end
		if(vga_x >= 10*width && vga_x < 11*width) begin
			background_x = 10*width;
			tile_x = 10;
		end
		if(vga_x >= 11*width && vga_x < 12*width) begin
			background_x = 11*width;
			tile_x = 11;
		end
		if(vga_x >= 12*width && vga_x < 13*width) begin
			background_x = 12*width;
			tile_x = 12;
		end
		if(vga_x >= 13*width && vga_x < 14*width) begin
			background_x = 13*width;
			tile_x = 13;
		end
		if(vga_x >= 14*width && vga_x < 15*width) begin
			background_x = 14*width;
			tile_x = 14;
		end
		if(vga_x >= 15*width && vga_x < 16*width) begin
			background_x = 15*width;
			tile_x = 15;
		end
		if(vga_x >= 16*width && vga_x < 17*width) begin
			background_x = 16*width;
			tile_x = 16;
		end
		if(vga_x >= 17*width && vga_x < 18*width) begin
			background_x = 17*width;
			tile_x = 17;
		end
		if(vga_x >= 18*width && vga_x < 19*width) begin
			background_x = 18*width;
			tile_x = 18;
		end
		if(vga_x >= 19*width && vga_x < 20*width) begin
			background_x = 19*width;
			tile_x = 19;
		end
		if(vga_x >= 20*width && vga_x < 21*width) begin
			background_x = 20*width;
			tile_x = 20;
		end
		if(vga_x >= 21*width && vga_x < 22*width) begin
			background_x = 21*width;
			tile_x = 21;
		end
		
		
		if(vga_y >= 0 && vga_y < height) begin
			background_y = 0;
			tile_y = 0;
		end
		if(vga_y >= height && vga_y < 2*height) begin
			background_y = height;
			tile_y = 1;
		end
		if(vga_y >= 2*height && vga_y < 3*height) begin
			background_y = 2*height;
			tile_y = 2;
		end
		if(vga_y >= 3*height && vga_y < 4*height) begin
			background_y = 3*height;
			tile_y = 3;
		end
		if(vga_y >= 4*height && vga_y < 5*height) begin
			background_y = 4*height;
			tile_y = 4;
		end
		if(vga_y >= 5*height && vga_y	< 6*height) begin
			background_y = 5*height;
			tile_y = 5;
		end
		if(vga_y >= 6*height && vga_y < 7*height) begin
			background_y = 6*height;
			tile_y = 6;
		end
		if(vga_y >= 7*height && vga_y < 8*height) begin
			background_y = 7*height;
			tile_y = 7;
		end
		if(vga_y >= 8*height && vga_y < 9*height) begin
			background_y = 8*height;
			tile_y = 8;
		end
		if(vga_y >= 9*height && vga_y < 10*height) begin
			background_y = 9*height;
			tile_y = 9;
		end
		if(vga_y >= 10*height && vga_y < 11*height) begin
			background_y = 10*height;
			tile_y = 10;
		end
		if(vga_y >= 11*height && vga_y < 12*height) begin
			background_y = 11*height;
			tile_y = 11;
		end
		if(vga_y >= 12*height && vga_y < 13*height) begin
			background_y = 12*height;
			tile_y = 12;
		end
		if(vga_y >= 13*height && vga_y < 14*height) begin
			background_y = 13*height;
			tile_y = 13;
		end
		if(vga_y >= 14*height && vga_y < 15*height) begin
			background_y = 14*height;
			tile_y = 14;
		end
		if(vga_y >= 15*height && vga_y < 16*height) begin
			background_y = 15*height;
			tile_y = 15;
		end
	end
	
	// Select the correct background tile from the background tile array:
	always_comb begin
		 // Default == Black
		 color = 33;
		 case(dummy[tile_y][tile_x])
			 0: begin
				color = BG1[vga_y - background_y][vga_x - background_x];
			 end
			 1: begin
				color = BG2[vga_y - background_y][vga_x - background_x];
			 end
			 2: begin
				color = BG3[vga_y - background_y][vga_x - background_x];
			 end
			 3: begin
				color = BG4[vga_y - background_y][vga_x - background_x];
			 end
			 4: begin
				color = BG5[vga_y - background_y][vga_x - background_x];
			 end
			 5: begin
				color = BG6[vga_y - background_y][vga_x - background_x];
			 end
			 6: begin
				color = BG7[vga_y - background_y][vga_x - background_x];
			 end
			 7: begin
				color = BG8[vga_y - background_y][vga_x - background_x];
			 end
			 default: begin
				color = 8;
			 end
		 endcase
		 if(color  == 0) color = 33;
	end
endmodule
